/******************************************************************************
 ** Logisim goes FPGA automatic generated Verilog code                       **
 **                                                                          **
 ** Component : RegFIle                                                      **
 **                                                                          **
 ******************************************************************************/

`timescale 1ns/1ps
module RegFIle( Clk,
                Din,
                LOGISIM_CLOCK_TREE_0,
                R1Adr,
                R2Adr,
                WAdr,
                WE,
                R1,
                R2);

   /***************************************************************************
    ** Here the inputs are defined                                           **
    ***************************************************************************/
   input  Clk;
   input[31:0]  Din;
   input[4:0]  LOGISIM_CLOCK_TREE_0;
   input[4:0]  R1Adr;
   input[4:0]  R2Adr;
   input[4:0]  WAdr;
   input  WE;

   /***************************************************************************
    ** Here the outputs are defined                                          **
    ***************************************************************************/
   output[31:0] R1;
   output[31:0] R2;

   /***************************************************************************
    ** Here the internal wires are defined                                   **
    ***************************************************************************/
   wire[31:0] s_LOGISIM_BUS_100;
   wire[31:0] s_LOGISIM_BUS_101;
   wire[31:0] s_LOGISIM_BUS_102;
   wire[31:0] s_LOGISIM_BUS_103;
   wire[31:0] s_LOGISIM_BUS_108;
   wire[31:0] s_LOGISIM_BUS_109;
   wire[31:0] s_LOGISIM_BUS_110;
   wire[31:0] s_LOGISIM_BUS_111;
   wire[31:0] s_LOGISIM_BUS_116;
   wire[31:0] s_LOGISIM_BUS_117;
   wire[31:0] s_LOGISIM_BUS_122;
   wire[31:0] s_LOGISIM_BUS_123;
   wire[31:0] s_LOGISIM_BUS_124;
   wire[31:0] s_LOGISIM_BUS_125;
   wire[31:0] s_LOGISIM_BUS_132;
   wire[31:0] s_LOGISIM_BUS_133;
   wire[31:0] s_LOGISIM_BUS_134;
   wire[31:0] s_LOGISIM_BUS_135;
   wire[31:0] s_LOGISIM_BUS_136;
   wire[31:0] s_LOGISIM_BUS_18;
   wire[4:0] s_LOGISIM_BUS_25;
   wire[4:0] s_LOGISIM_BUS_26;
   wire[31:0] s_LOGISIM_BUS_36;
   wire[31:0] s_LOGISIM_BUS_37;
   wire[31:0] s_LOGISIM_BUS_46;
   wire[31:0] s_LOGISIM_BUS_48;
   wire[31:0] s_LOGISIM_BUS_56;
   wire[31:0] s_LOGISIM_BUS_57;
   wire[31:0] s_LOGISIM_BUS_6;
   wire[31:0] s_LOGISIM_BUS_66;
   wire[31:0] s_LOGISIM_BUS_67;
   wire[31:0] s_LOGISIM_BUS_75;
   wire[31:0] s_LOGISIM_BUS_76;
   wire[31:0] s_LOGISIM_BUS_85;
   wire[31:0] s_LOGISIM_BUS_86;
   wire[31:0] s_LOGISIM_BUS_87;
   wire[31:0] s_LOGISIM_BUS_88;
   wire[31:0] s_LOGISIM_BUS_94;
   wire[4:0] s_LOGISIM_BUS_97;
   wire s_LOGISIM_NET_0;
   wire s_LOGISIM_NET_1;
   wire s_LOGISIM_NET_10;
   wire s_LOGISIM_NET_104;
   wire s_LOGISIM_NET_105;
   wire s_LOGISIM_NET_106;
   wire s_LOGISIM_NET_107;
   wire s_LOGISIM_NET_11;
   wire s_LOGISIM_NET_112;
   wire s_LOGISIM_NET_113;
   wire s_LOGISIM_NET_114;
   wire s_LOGISIM_NET_115;
   wire s_LOGISIM_NET_118;
   wire s_LOGISIM_NET_119;
   wire s_LOGISIM_NET_12;
   wire s_LOGISIM_NET_120;
   wire s_LOGISIM_NET_121;
   wire s_LOGISIM_NET_126;
   wire s_LOGISIM_NET_127;
   wire s_LOGISIM_NET_128;
   wire s_LOGISIM_NET_129;
   wire s_LOGISIM_NET_13;
   wire s_LOGISIM_NET_130;
   wire s_LOGISIM_NET_131;
   wire s_LOGISIM_NET_137;
   wire s_LOGISIM_NET_138;
   wire s_LOGISIM_NET_139;
   wire s_LOGISIM_NET_14;
   wire s_LOGISIM_NET_140;
   wire s_LOGISIM_NET_141;
   wire s_LOGISIM_NET_142;
   wire s_LOGISIM_NET_143;
   wire s_LOGISIM_NET_144;
   wire s_LOGISIM_NET_145;
   wire s_LOGISIM_NET_146;
   wire s_LOGISIM_NET_147;
   wire s_LOGISIM_NET_148;
   wire s_LOGISIM_NET_149;
   wire s_LOGISIM_NET_15;
   wire s_LOGISIM_NET_150;
   wire s_LOGISIM_NET_151;
   wire s_LOGISIM_NET_152;
   wire s_LOGISIM_NET_153;
   wire s_LOGISIM_NET_154;
   wire s_LOGISIM_NET_155;
   wire s_LOGISIM_NET_156;
   wire s_LOGISIM_NET_157;
   wire s_LOGISIM_NET_158;
   wire s_LOGISIM_NET_159;
   wire s_LOGISIM_NET_16;
   wire s_LOGISIM_NET_160;
   wire s_LOGISIM_NET_161;
   wire s_LOGISIM_NET_162;
   wire s_LOGISIM_NET_163;
   wire s_LOGISIM_NET_164;
   wire s_LOGISIM_NET_165;
   wire s_LOGISIM_NET_166;
   wire s_LOGISIM_NET_167;
   wire s_LOGISIM_NET_168;
   wire s_LOGISIM_NET_17;
   wire s_LOGISIM_NET_19;
   wire s_LOGISIM_NET_2;
   wire s_LOGISIM_NET_20;
   wire s_LOGISIM_NET_21;
   wire s_LOGISIM_NET_22;
   wire s_LOGISIM_NET_23;
   wire s_LOGISIM_NET_24;
   wire s_LOGISIM_NET_27;
   wire s_LOGISIM_NET_28;
   wire s_LOGISIM_NET_29;
   wire s_LOGISIM_NET_3;
   wire s_LOGISIM_NET_30;
   wire s_LOGISIM_NET_31;
   wire s_LOGISIM_NET_32;
   wire s_LOGISIM_NET_33;
   wire s_LOGISIM_NET_34;
   wire s_LOGISIM_NET_35;
   wire s_LOGISIM_NET_38;
   wire s_LOGISIM_NET_39;
   wire s_LOGISIM_NET_4;
   wire s_LOGISIM_NET_40;
   wire s_LOGISIM_NET_41;
   wire s_LOGISIM_NET_42;
   wire s_LOGISIM_NET_43;
   wire s_LOGISIM_NET_44;
   wire s_LOGISIM_NET_45;
   wire s_LOGISIM_NET_47;
   wire s_LOGISIM_NET_49;
   wire s_LOGISIM_NET_5;
   wire s_LOGISIM_NET_50;
   wire s_LOGISIM_NET_51;
   wire s_LOGISIM_NET_52;
   wire s_LOGISIM_NET_53;
   wire s_LOGISIM_NET_54;
   wire s_LOGISIM_NET_55;
   wire s_LOGISIM_NET_58;
   wire s_LOGISIM_NET_59;
   wire s_LOGISIM_NET_60;
   wire s_LOGISIM_NET_61;
   wire s_LOGISIM_NET_62;
   wire s_LOGISIM_NET_63;
   wire s_LOGISIM_NET_64;
   wire s_LOGISIM_NET_65;
   wire s_LOGISIM_NET_68;
   wire s_LOGISIM_NET_69;
   wire s_LOGISIM_NET_7;
   wire s_LOGISIM_NET_70;
   wire s_LOGISIM_NET_71;
   wire s_LOGISIM_NET_72;
   wire s_LOGISIM_NET_73;
   wire s_LOGISIM_NET_74;
   wire s_LOGISIM_NET_77;
   wire s_LOGISIM_NET_78;
   wire s_LOGISIM_NET_79;
   wire s_LOGISIM_NET_8;
   wire s_LOGISIM_NET_80;
   wire s_LOGISIM_NET_81;
   wire s_LOGISIM_NET_82;
   wire s_LOGISIM_NET_83;
   wire s_LOGISIM_NET_84;
   wire s_LOGISIM_NET_89;
   wire s_LOGISIM_NET_9;
   wire s_LOGISIM_NET_90;
   wire s_LOGISIM_NET_91;
   wire s_LOGISIM_NET_92;
   wire s_LOGISIM_NET_93;
   wire s_LOGISIM_NET_95;
   wire s_LOGISIM_NET_96;
   wire s_LOGISIM_NET_98;
   wire s_LOGISIM_NET_99;


   /***************************************************************************
    ** Here all input connections are defined                                **
    ***************************************************************************/
   assign s_LOGISIM_BUS_136[31:0]            = Din;
   assign s_LOGISIM_NET_38                   = WE;
   assign s_LOGISIM_BUS_97[4:0]              = WAdr;
   assign s_LOGISIM_NET_131                  = Clk;
   assign s_LOGISIM_BUS_26[4:0]              = R2Adr;
   assign s_LOGISIM_BUS_25[4:0]              = R1Adr;

   /***************************************************************************
    ** Here all output connections are defined                               **
    ***************************************************************************/
   assign R1                                 = s_LOGISIM_BUS_46[31:0];
   assign R2                                 = s_LOGISIM_BUS_6[31:0];

   /***************************************************************************
    ** Here all in-lined components are defined                              **
    ***************************************************************************/
   assign s_LOGISIM_NET_8 = 1'd0;

   assign s_LOGISIM_NET_165 = 1'd0;

   assign s_LOGISIM_NET_141 = 1'd0;

   assign s_LOGISIM_NET_53 = 1'd0;

   assign s_LOGISIM_NET_128 = 1'd0;

   assign s_LOGISIM_NET_49 = 1'd0;

   assign s_LOGISIM_NET_164 = 1'd0;

   assign s_LOGISIM_NET_161 = 1'd0;

   assign s_LOGISIM_NET_50 = 1'd0;

   assign s_LOGISIM_NET_106 = 1'd0;

   assign s_LOGISIM_BUS_103[31:0] = 32'd0;

   assign s_LOGISIM_NET_140 = 1'd0;

   assign s_LOGISIM_NET_5 = 1'd0;

   assign s_LOGISIM_NET_0 = 1'd0;

   assign s_LOGISIM_NET_148 = 1'd0;

   assign s_LOGISIM_NET_163 = 1'd0;

   assign s_LOGISIM_NET_42 = 1'd0;

   assign s_LOGISIM_NET_167 = 1'd0;

   assign s_LOGISIM_NET_9 = 1'd0;

   assign s_LOGISIM_NET_74 = 1'd0;

   assign s_LOGISIM_NET_142 = 1'd0;

   assign s_LOGISIM_NET_52 = 1'd0;

   assign s_LOGISIM_NET_146 = 1'd0;

   assign s_LOGISIM_NET_143 = 1'd0;

   assign s_LOGISIM_NET_40 = 1'd0;

   assign s_LOGISIM_NET_62 = 1'd0;

   assign s_LOGISIM_NET_61 = 1'd0;

   assign s_LOGISIM_NET_153 = 1'd0;

   assign s_LOGISIM_NET_33 = 1'd0;

   assign s_LOGISIM_NET_44 = 1'd0;

   assign s_LOGISIM_NET_139 = 1'd0;

   assign s_LOGISIM_NET_145 = 1'd0;

   assign s_LOGISIM_NET_21 = 1'd0;

   assign s_LOGISIM_NET_14 = 1'd0;

   assign s_LOGISIM_NET_19 = 1'd0;

   assign s_LOGISIM_NET_32 = 1'd0;

   assign s_LOGISIM_NET_72 = 1'd0;

   assign s_LOGISIM_NET_81 = 1'd0;

   assign s_LOGISIM_NET_144 = 1'd0;

   assign s_LOGISIM_NET_45 = 1'd0;

   assign s_LOGISIM_NET_126 = 1'd0;

   assign s_LOGISIM_NET_20 = 1'd0;

   assign s_LOGISIM_NET_35 = 1'd0;

   assign s_LOGISIM_NET_17 = 1'd0;

   assign s_LOGISIM_NET_54 = 1'd0;

   assign s_LOGISIM_NET_149 = 1'd0;

   assign s_LOGISIM_NET_2 = 1'd0;

   assign s_LOGISIM_NET_121 = 1'd0;

   assign s_LOGISIM_NET_147 = 1'd0;

   assign s_LOGISIM_NET_1 = 1'd0;

   assign s_LOGISIM_NET_3 = 1'd0;

   assign s_LOGISIM_NET_4 = 1'd0;

   assign s_LOGISIM_NET_118 = 1'd0;

   assign s_LOGISIM_NET_150 = 1'd0;

   assign s_LOGISIM_NET_151 = 1'd0;

   assign s_LOGISIM_NET_43 = 1'd0;

   assign s_LOGISIM_NET_15 = 1'd0;

   assign s_LOGISIM_NET_68 = 1'd0;

   assign s_LOGISIM_NET_27 = 1'd0;

   assign s_LOGISIM_NET_113 = 1'd0;

   assign s_LOGISIM_NET_12 = 1'd0;

   assign s_LOGISIM_NET_152 = 1'd0;

   assign s_LOGISIM_NET_7 = 1'd0;

   assign s_LOGISIM_NET_154 = 1'd0;

   assign s_LOGISIM_NET_155 = 1'd0;

   assign s_LOGISIM_NET_156 = 1'd0;

   assign s_LOGISIM_NET_24 = 1'd0;

   assign s_LOGISIM_NET_91 = 1'd0;

   assign s_LOGISIM_NET_78 = 1'd0;

   assign s_LOGISIM_NET_127 = 1'd0;

   assign s_LOGISIM_NET_23 = 1'd0;

   assign s_LOGISIM_NET_34 = 1'd0;

   assign s_LOGISIM_NET_157 = 1'd0;

   assign s_LOGISIM_NET_158 = 1'd0;

   assign s_LOGISIM_NET_10 = 1'd0;

   assign s_LOGISIM_NET_159 = 1'd0;

   assign s_LOGISIM_NET_160 = 1'd0;

   assign s_LOGISIM_NET_95 = 1'd0;

   assign s_LOGISIM_NET_22 = 1'd0;

   assign s_LOGISIM_NET_162 = 1'd0;

   assign s_LOGISIM_NET_69 = 1'd0;

   assign s_LOGISIM_NET_63 = 1'd0;

   assign s_LOGISIM_NET_112 = 1'd0;

   assign s_LOGISIM_NET_47 = 1'd0;

   assign s_LOGISIM_NET_166 = 1'd0;

   assign s_LOGISIM_NET_13 = 1'd0;

   assign s_LOGISIM_NET_93 = 1'd0;

   assign s_LOGISIM_NET_41 = 1'd0;

   assign s_LOGISIM_NET_59 = 1'd0;

   assign s_LOGISIM_NET_96 = 1'd0;

   assign s_LOGISIM_NET_82 = 1'd0;

   assign s_LOGISIM_NET_16 = 1'd0;

   assign s_LOGISIM_NET_55 = 1'd0;

   assign s_LOGISIM_NET_80 = 1'd0;

   assign s_LOGISIM_NET_168 = 1'd0;

   assign s_LOGISIM_NET_28 = 1'd0;

   assign s_LOGISIM_NET_107 = 1'd0;


   /***************************************************************************
    ** Here all normal components are defined                                **
    ***************************************************************************/
   REGISTER_FLIP_FLOP_s28 #(.ActiveLevel(1),
                            .NrOfBits(32))
      REGISTER_FILE_1 (.Clock(LOGISIM_CLOCK_TREE_0[4]),
                       .ClockEnable(s_LOGISIM_NET_90),
                       .D(s_LOGISIM_BUS_136[31:0]),
                       .Q(s_LOGISIM_BUS_102[31:0]),
                       .Reset(s_LOGISIM_NET_9),
                       .Tick(LOGISIM_CLOCK_TREE_0[2]),
                       .cs(s_LOGISIM_NET_52),
                       .pre(s_LOGISIM_NET_143));

   REGISTER_FLIP_FLOP_s21 #(.ActiveLevel(1),
                            .NrOfBits(32))
      REGISTER_FILE_2 (.Clock(LOGISIM_CLOCK_TREE_0[4]),
                       .ClockEnable(s_LOGISIM_NET_130),
                       .D(s_LOGISIM_BUS_136[31:0]),
                       .Q(s_LOGISIM_BUS_116[31:0]),
                       .Reset(s_LOGISIM_NET_24),
                       .Tick(LOGISIM_CLOCK_TREE_0[2]),
                       .cs(s_LOGISIM_NET_74),
                       .pre(s_LOGISIM_NET_147));

   REGISTER_FLIP_FLOP_s9 #(.ActiveLevel(1),
                           .NrOfBits(32))
      REGISTER_FILE_3 (.Clock(LOGISIM_CLOCK_TREE_0[4]),
                       .ClockEnable(s_LOGISIM_NET_77),
                       .D(s_LOGISIM_BUS_136[31:0]),
                       .Q(s_LOGISIM_BUS_122[31:0]),
                       .Reset(s_LOGISIM_NET_3),
                       .Tick(LOGISIM_CLOCK_TREE_0[2]),
                       .cs(s_LOGISIM_NET_40),
                       .pre(s_LOGISIM_NET_141));

   REGISTER_FLIP_FLOP_s16 #(.ActiveLevel(1),
                            .NrOfBits(32))
      REGISTER_FILE_4 (.Clock(LOGISIM_CLOCK_TREE_0[4]),
                       .ClockEnable(s_LOGISIM_NET_120),
                       .D(s_LOGISIM_BUS_136[31:0]),
                       .Q(s_LOGISIM_BUS_134[31:0]),
                       .Reset(s_LOGISIM_NET_22),
                       .Tick(LOGISIM_CLOCK_TREE_0[2]),
                       .cs(s_LOGISIM_NET_118),
                       .pre(s_LOGISIM_NET_1));

   REGISTER_FLIP_FLOP_s2 #(.ActiveLevel(1),
                           .NrOfBits(32))
      REGISTER_FILE_5 (.Clock(LOGISIM_CLOCK_TREE_0[4]),
                       .ClockEnable(s_LOGISIM_NET_70),
                       .D(s_LOGISIM_BUS_136[31:0]),
                       .Q(s_LOGISIM_BUS_88[31:0]),
                       .Reset(s_LOGISIM_NET_50),
                       .Tick(LOGISIM_CLOCK_TREE_0[2]),
                       .cs(s_LOGISIM_NET_5),
                       .pre(s_LOGISIM_NET_154));

   REGISTER_FLIP_FLOP_s24 #(.ActiveLevel(1),
                            .NrOfBits(32))
      REGISTER_FILE_6 (.Clock(LOGISIM_CLOCK_TREE_0[4]),
                       .ClockEnable(s_LOGISIM_NET_51),
                       .D(s_LOGISIM_BUS_136[31:0]),
                       .Q(s_LOGISIM_BUS_67[31:0]),
                       .Reset(s_LOGISIM_NET_21),
                       .Tick(LOGISIM_CLOCK_TREE_0[2]),
                       .cs(s_LOGISIM_NET_121),
                       .pre(s_LOGISIM_NET_0));

   REGISTER_FLIP_FLOP_s5 #(.ActiveLevel(1),
                           .NrOfBits(32))
      REGISTER_FILE_7 (.Clock(LOGISIM_CLOCK_TREE_0[4]),
                       .ClockEnable(s_LOGISIM_NET_129),
                       .D(s_LOGISIM_BUS_136[31:0]),
                       .Q(s_LOGISIM_BUS_111[31:0]),
                       .Reset(s_LOGISIM_NET_16),
                       .Tick(LOGISIM_CLOCK_TREE_0[2]),
                       .cs(s_LOGISIM_NET_61),
                       .pre(s_LOGISIM_NET_159));

   REGISTER_FLIP_FLOP_s31 #(.ActiveLevel(1),
                            .NrOfBits(32))
      REGISTER_FILE_8 (.Clock(LOGISIM_CLOCK_TREE_0[4]),
                       .ClockEnable(s_LOGISIM_NET_11),
                       .D(s_LOGISIM_BUS_136[31:0]),
                       .Q(s_LOGISIM_BUS_109[31:0]),
                       .Reset(s_LOGISIM_NET_7),
                       .Tick(LOGISIM_CLOCK_TREE_0[2]),
                       .cs(s_LOGISIM_NET_106),
                       .pre(s_LOGISIM_NET_162));

   REGISTER_FLIP_FLOP_s15 #(.ActiveLevel(1),
                            .NrOfBits(32))
      REGISTER_FILE_9 (.Clock(LOGISIM_CLOCK_TREE_0[4]),
                       .ClockEnable(s_LOGISIM_NET_39),
                       .D(s_LOGISIM_BUS_136[31:0]),
                       .Q(s_LOGISIM_BUS_108[31:0]),
                       .Reset(s_LOGISIM_NET_49),
                       .Tick(LOGISIM_CLOCK_TREE_0[2]),
                       .cs(s_LOGISIM_NET_4),
                       .pre(s_LOGISIM_NET_152));

   REGISTER_FLIP_FLOP_s14 #(.ActiveLevel(1),
                            .NrOfBits(32))
      REGISTER_FILE_10 (.Clock(LOGISIM_CLOCK_TREE_0[4]),
                        .ClockEnable(s_LOGISIM_NET_29),
                        .D(s_LOGISIM_BUS_136[31:0]),
                        .Q(s_LOGISIM_BUS_48[31:0]),
                        .Reset(s_LOGISIM_NET_27),
                        .Tick(LOGISIM_CLOCK_TREE_0[2]),
                        .cs(s_LOGISIM_NET_126),
                        .pre(s_LOGISIM_NET_142));

   REGISTER_FLIP_FLOP_s18 #(.ActiveLevel(1),
                            .NrOfBits(32))
      REGISTER_FILE_11 (.Clock(LOGISIM_CLOCK_TREE_0[4]),
                        .ClockEnable(s_LOGISIM_NET_71),
                        .D(s_LOGISIM_BUS_136[31:0]),
                        .Q(s_LOGISIM_BUS_87[31:0]),
                        .Reset(s_LOGISIM_NET_63),
                        .Tick(LOGISIM_CLOCK_TREE_0[2]),
                        .cs(s_LOGISIM_NET_15),
                        .pre(s_LOGISIM_NET_155));

   REGISTER_FLIP_FLOP_s8 #(.ActiveLevel(1),
                           .NrOfBits(32))
      REGISTER_FILE_12 (.Clock(LOGISIM_CLOCK_TREE_0[4]),
                        .ClockEnable(s_LOGISIM_NET_58),
                        .D(s_LOGISIM_BUS_136[31:0]),
                        .Q(s_LOGISIM_BUS_75[31:0]),
                        .Reset(s_LOGISIM_NET_68),
                        .Tick(LOGISIM_CLOCK_TREE_0[2]),
                        .cs(s_LOGISIM_NET_19),
                        .pre(s_LOGISIM_NET_47));

   REGISTER_FLIP_FLOP_s19 #(.ActiveLevel(1),
                            .NrOfBits(32))
      REGISTER_FILE_13 (.Clock(LOGISIM_CLOCK_TREE_0[4]),
                        .ClockEnable(s_LOGISIM_NET_73),
                        .D(s_LOGISIM_BUS_136[31:0]),
                        .Q(s_LOGISIM_BUS_85[31:0]),
                        .Reset(s_LOGISIM_NET_82),
                        .Tick(LOGISIM_CLOCK_TREE_0[2]),
                        .cs(s_LOGISIM_NET_33),
                        .pre(s_LOGISIM_NET_151));

   REGISTER_FLIP_FLOP_s10 #(.ActiveLevel(1),
                            .NrOfBits(32))
      REGISTER_FILE_14 (.Clock(LOGISIM_CLOCK_TREE_0[4]),
                        .ClockEnable(s_LOGISIM_NET_137),
                        .D(s_LOGISIM_BUS_136[31:0]),
                        .Q(s_LOGISIM_BUS_110[31:0]),
                        .Reset(s_LOGISIM_NET_17),
                        .Tick(LOGISIM_CLOCK_TREE_0[2]),
                        .cs(s_LOGISIM_NET_59),
                        .pre(s_LOGISIM_NET_144));

   REGISTER_FLIP_FLOP_s20 #(.ActiveLevel(1),
                            .NrOfBits(32))
      REGISTER_FILE_15 (.Clock(LOGISIM_CLOCK_TREE_0[4]),
                        .ClockEnable(s_LOGISIM_NET_92),
                        .D(s_LOGISIM_BUS_136[31:0]),
                        .Q(s_LOGISIM_BUS_100[31:0]),
                        .Reset(s_LOGISIM_NET_10),
                        .Tick(LOGISIM_CLOCK_TREE_0[2]),
                        .cs(s_LOGISIM_NET_53),
                        .pre(s_LOGISIM_NET_157));

   REGISTER_FLIP_FLOP_s25 #(.ActiveLevel(1),
                            .NrOfBits(32))
      REGISTER_FILE_16 (.Clock(LOGISIM_CLOCK_TREE_0[4]),
                        .ClockEnable(s_LOGISIM_NET_31),
                        .D(s_LOGISIM_BUS_136[31:0]),
                        .Q(s_LOGISIM_BUS_123[31:0]),
                        .Reset(s_LOGISIM_NET_42),
                        .Tick(LOGISIM_CLOCK_TREE_0[2]),
                        .cs(s_LOGISIM_NET_139),
                        .pre(s_LOGISIM_NET_145));

   REGISTER_FLIP_FLOP_s3 #(.ActiveLevel(1),
                           .NrOfBits(32))
      REGISTER_FILE_17 (.Clock(LOGISIM_CLOCK_TREE_0[4]),
                        .ClockEnable(s_LOGISIM_NET_60),
                        .D(s_LOGISIM_BUS_136[31:0]),
                        .Q(s_LOGISIM_BUS_76[31:0]),
                        .Reset(s_LOGISIM_NET_69),
                        .Tick(LOGISIM_CLOCK_TREE_0[2]),
                        .cs(s_LOGISIM_NET_20),
                        .pre(s_LOGISIM_NET_146));

   REGISTER_FLIP_FLOP_s30 #(.ActiveLevel(1),
                            .NrOfBits(32))
      REGISTER_FILE_18 (.Clock(LOGISIM_CLOCK_TREE_0[4]),
                        .ClockEnable(s_LOGISIM_NET_30),
                        .D(s_LOGISIM_BUS_136[31:0]),
                        .Q(s_LOGISIM_BUS_133[31:0]),
                        .Reset(s_LOGISIM_NET_44),
                        .Tick(LOGISIM_CLOCK_TREE_0[2]),
                        .cs(s_LOGISIM_NET_91),
                        .pre(s_LOGISIM_NET_166));

   REGISTER_FLIP_FLOP_s17 #(.ActiveLevel(1),
                            .NrOfBits(32))
      REGISTER_FILE_19 (.Clock(LOGISIM_CLOCK_TREE_0[4]),
                        .ClockEnable(s_LOGISIM_NET_99),
                        .D(s_LOGISIM_BUS_136[31:0]),
                        .Q(s_LOGISIM_BUS_57[31:0]),
                        .Reset(s_LOGISIM_NET_43),
                        .Tick(LOGISIM_CLOCK_TREE_0[2]),
                        .cs(s_LOGISIM_NET_140),
                        .pre(s_LOGISIM_NET_148));

   REGISTER_FLIP_FLOP_s29 #(.ActiveLevel(1),
                            .NrOfBits(32))
      REGISTER_FILE_20 (.Clock(LOGISIM_CLOCK_TREE_0[4]),
                        .ClockEnable(s_LOGISIM_NET_65),
                        .D(s_LOGISIM_BUS_136[31:0]),
                        .Q(s_LOGISIM_BUS_117[31:0]),
                        .Reset(s_LOGISIM_NET_23),
                        .Tick(LOGISIM_CLOCK_TREE_0[2]),
                        .cs(s_LOGISIM_NET_72),
                        .pre(s_LOGISIM_NET_149));

   REGISTER_FLIP_FLOP_s26 #(.ActiveLevel(1),
                            .NrOfBits(32))
      REGISTER_FILE_21 (.Clock(LOGISIM_CLOCK_TREE_0[4]),
                        .ClockEnable(s_LOGISIM_NET_138),
                        .D(s_LOGISIM_BUS_136[31:0]),
                        .Q(s_LOGISIM_BUS_66[31:0]),
                        .Reset(s_LOGISIM_NET_62),
                        .Tick(LOGISIM_CLOCK_TREE_0[2]),
                        .cs(s_LOGISIM_NET_14),
                        .pre(s_LOGISIM_NET_150));

   Demultiplexer_32      DEMUX_1 (.DemuxIn(s_LOGISIM_NET_38),
                                  .DemuxOut_0(s_LOGISIM_NET_119),
                                  .DemuxOut_1(s_LOGISIM_NET_98),
                                  .DemuxOut_10(s_LOGISIM_NET_137),
                                  .DemuxOut_11(s_LOGISIM_NET_114),
                                  .DemuxOut_12(s_LOGISIM_NET_89),
                                  .DemuxOut_13(s_LOGISIM_NET_64),
                                  .DemuxOut_14(s_LOGISIM_NET_29),
                                  .DemuxOut_15(s_LOGISIM_NET_39),
                                  .DemuxOut_16(s_LOGISIM_NET_120),
                                  .DemuxOut_17(s_LOGISIM_NET_99),
                                  .DemuxOut_18(s_LOGISIM_NET_71),
                                  .DemuxOut_19(s_LOGISIM_NET_73),
                                  .DemuxOut_2(s_LOGISIM_NET_70),
                                  .DemuxOut_20(s_LOGISIM_NET_92),
                                  .DemuxOut_21(s_LOGISIM_NET_130),
                                  .DemuxOut_22(s_LOGISIM_NET_105),
                                  .DemuxOut_23(s_LOGISIM_NET_84),
                                  .DemuxOut_24(s_LOGISIM_NET_51),
                                  .DemuxOut_25(s_LOGISIM_NET_31),
                                  .DemuxOut_26(s_LOGISIM_NET_138),
                                  .DemuxOut_27(s_LOGISIM_NET_115),
                                  .DemuxOut_28(s_LOGISIM_NET_90),
                                  .DemuxOut_29(s_LOGISIM_NET_65),
                                  .DemuxOut_3(s_LOGISIM_NET_60),
                                  .DemuxOut_30(s_LOGISIM_NET_30),
                                  .DemuxOut_31(s_LOGISIM_NET_11),
                                  .DemuxOut_4(s_LOGISIM_NET_79),
                                  .DemuxOut_5(s_LOGISIM_NET_129),
                                  .DemuxOut_6(s_LOGISIM_NET_104),
                                  .DemuxOut_7(s_LOGISIM_NET_83),
                                  .DemuxOut_8(s_LOGISIM_NET_58),
                                  .DemuxOut_9(s_LOGISIM_NET_77),
                                  .Enable(1'b1),
                                  .Sel(s_LOGISIM_BUS_97[4:0]));

   REGISTER_FLIP_FLOP_s13 #(.ActiveLevel(1),
                            .NrOfBits(32))
      REGISTER_FILE_22 (.Clock(LOGISIM_CLOCK_TREE_0[4]),
                        .ClockEnable(s_LOGISIM_NET_64),
                        .D(s_LOGISIM_BUS_136[31:0]),
                        .Q(s_LOGISIM_BUS_18[31:0]),
                        .Reset(s_LOGISIM_NET_12),
                        .Tick(LOGISIM_CLOCK_TREE_0[2]),
                        .cs(s_LOGISIM_NET_112),
                        .pre(s_LOGISIM_NET_153));

   REGISTER_FLIP_FLOP_s27 #(.ActiveLevel(1),
                            .NrOfBits(32))
      REGISTER_FILE_23 (.Clock(LOGISIM_CLOCK_TREE_0[4]),
                        .ClockEnable(s_LOGISIM_NET_115),
                        .D(s_LOGISIM_BUS_136[31:0]),
                        .Q(s_LOGISIM_BUS_86[31:0]),
                        .Reset(s_LOGISIM_NET_81),
                        .Tick(LOGISIM_CLOCK_TREE_0[2]),
                        .cs(s_LOGISIM_NET_32),
                        .pre(s_LOGISIM_NET_156));

   REGISTER_FLIP_FLOP_s11 #(.ActiveLevel(1),
                            .NrOfBits(32))
      REGISTER_FILE_24 (.Clock(LOGISIM_CLOCK_TREE_0[4]),
                        .ClockEnable(s_LOGISIM_NET_114),
                        .D(s_LOGISIM_BUS_136[31:0]),
                        .Q(s_LOGISIM_BUS_124[31:0]),
                        .Reset(s_LOGISIM_NET_35),
                        .Tick(LOGISIM_CLOCK_TREE_0[2]),
                        .cs(s_LOGISIM_NET_78),
                        .pre(s_LOGISIM_NET_158));

   REGISTER_FLIP_FLOP_s1 #(.ActiveLevel(1),
                           .NrOfBits(32))
      REGISTER_FILE_25 (.Clock(LOGISIM_CLOCK_TREE_0[4]),
                        .ClockEnable(s_LOGISIM_NET_98),
                        .D(s_LOGISIM_BUS_136[31:0]),
                        .Q(s_LOGISIM_BUS_56[31:0]),
                        .Reset(s_LOGISIM_NET_28),
                        .Tick(LOGISIM_CLOCK_TREE_0[2]),
                        .cs(s_LOGISIM_NET_127),
                        .pre(s_LOGISIM_NET_160));

   REGISTER_FLIP_FLOP_s23 #(.ActiveLevel(1),
                            .NrOfBits(32))
      REGISTER_FILE_26 (.Clock(LOGISIM_CLOCK_TREE_0[4]),
                        .ClockEnable(s_LOGISIM_NET_84),
                        .D(s_LOGISIM_BUS_136[31:0]),
                        .Q(s_LOGISIM_BUS_37[31:0]),
                        .Reset(s_LOGISIM_NET_8),
                        .Tick(LOGISIM_CLOCK_TREE_0[2]),
                        .cs(s_LOGISIM_NET_107),
                        .pre(s_LOGISIM_NET_161));

   REGISTER_FLIP_FLOP_s0 #(.ActiveLevel(1),
                           .NrOfBits(32))
      REGISTER_FILE_27 (.Clock(LOGISIM_CLOCK_TREE_0[4]),
                        .ClockEnable(s_LOGISIM_NET_119),
                        .D(s_LOGISIM_BUS_103[31:0]),
                        .Q(s_LOGISIM_BUS_135[31:0]),
                        .Reset(s_LOGISIM_NET_13),
                        .Tick(LOGISIM_CLOCK_TREE_0[2]),
                        .cs(s_LOGISIM_NET_113),
                        .pre(s_LOGISIM_NET_128));

   REGISTER_FLIP_FLOP_s4 #(.ActiveLevel(1),
                           .NrOfBits(32))
      REGISTER_FILE_28 (.Clock(LOGISIM_CLOCK_TREE_0[4]),
                        .ClockEnable(s_LOGISIM_NET_79),
                        .D(s_LOGISIM_BUS_136[31:0]),
                        .Q(s_LOGISIM_BUS_94[31:0]),
                        .Reset(s_LOGISIM_NET_2),
                        .Tick(LOGISIM_CLOCK_TREE_0[2]),
                        .cs(s_LOGISIM_NET_41),
                        .pre(s_LOGISIM_NET_163));

   REGISTER_FLIP_FLOP_s7 #(.ActiveLevel(1),
                           .NrOfBits(32))
      REGISTER_FILE_29 (.Clock(LOGISIM_CLOCK_TREE_0[4]),
                        .ClockEnable(s_LOGISIM_NET_83),
                        .D(s_LOGISIM_BUS_136[31:0]),
                        .Q(s_LOGISIM_BUS_36[31:0]),
                        .Reset(s_LOGISIM_NET_54),
                        .Tick(LOGISIM_CLOCK_TREE_0[2]),
                        .cs(s_LOGISIM_NET_96),
                        .pre(s_LOGISIM_NET_164));

   REGISTER_FLIP_FLOP_s12 #(.ActiveLevel(1),
                            .NrOfBits(32))
      REGISTER_FILE_30 (.Clock(LOGISIM_CLOCK_TREE_0[4]),
                        .ClockEnable(s_LOGISIM_NET_89),
                        .D(s_LOGISIM_BUS_136[31:0]),
                        .Q(s_LOGISIM_BUS_101[31:0]),
                        .Reset(s_LOGISIM_NET_55),
                        .Tick(LOGISIM_CLOCK_TREE_0[2]),
                        .cs(s_LOGISIM_NET_95),
                        .pre(s_LOGISIM_NET_165));

   Multiplexer_bus_32 #(.NrOfBits(32))
      MUX_1 (.Enable(1'b1),
             .MuxIn_0(s_LOGISIM_BUS_135[31:0]),
             .MuxIn_1(s_LOGISIM_BUS_56[31:0]),
             .MuxIn_10(s_LOGISIM_BUS_110[31:0]),
             .MuxIn_11(s_LOGISIM_BUS_124[31:0]),
             .MuxIn_12(s_LOGISIM_BUS_101[31:0]),
             .MuxIn_13(s_LOGISIM_BUS_18[31:0]),
             .MuxIn_14(s_LOGISIM_BUS_48[31:0]),
             .MuxIn_15(s_LOGISIM_BUS_108[31:0]),
             .MuxIn_16(s_LOGISIM_BUS_134[31:0]),
             .MuxIn_17(s_LOGISIM_BUS_57[31:0]),
             .MuxIn_18(s_LOGISIM_BUS_87[31:0]),
             .MuxIn_19(s_LOGISIM_BUS_85[31:0]),
             .MuxIn_2(s_LOGISIM_BUS_88[31:0]),
             .MuxIn_20(s_LOGISIM_BUS_100[31:0]),
             .MuxIn_21(s_LOGISIM_BUS_116[31:0]),
             .MuxIn_22(s_LOGISIM_BUS_132[31:0]),
             .MuxIn_23(s_LOGISIM_BUS_37[31:0]),
             .MuxIn_24(s_LOGISIM_BUS_67[31:0]),
             .MuxIn_25(s_LOGISIM_BUS_123[31:0]),
             .MuxIn_26(s_LOGISIM_BUS_66[31:0]),
             .MuxIn_27(s_LOGISIM_BUS_86[31:0]),
             .MuxIn_28(s_LOGISIM_BUS_102[31:0]),
             .MuxIn_29(s_LOGISIM_BUS_117[31:0]),
             .MuxIn_3(s_LOGISIM_BUS_76[31:0]),
             .MuxIn_30(s_LOGISIM_BUS_133[31:0]),
             .MuxIn_31(s_LOGISIM_BUS_109[31:0]),
             .MuxIn_4(s_LOGISIM_BUS_94[31:0]),
             .MuxIn_5(s_LOGISIM_BUS_111[31:0]),
             .MuxIn_6(s_LOGISIM_BUS_125[31:0]),
             .MuxIn_7(s_LOGISIM_BUS_36[31:0]),
             .MuxIn_8(s_LOGISIM_BUS_75[31:0]),
             .MuxIn_9(s_LOGISIM_BUS_122[31:0]),
             .MuxOut(s_LOGISIM_BUS_46[31:0]),
             .Sel(s_LOGISIM_BUS_25[4:0]));

   REGISTER_FLIP_FLOP_s22 #(.ActiveLevel(1),
                            .NrOfBits(32))
      REGISTER_FILE_31 (.Clock(LOGISIM_CLOCK_TREE_0[4]),
                        .ClockEnable(s_LOGISIM_NET_105),
                        .D(s_LOGISIM_BUS_136[31:0]),
                        .Q(s_LOGISIM_BUS_132[31:0]),
                        .Reset(s_LOGISIM_NET_45),
                        .Tick(LOGISIM_CLOCK_TREE_0[2]),
                        .cs(s_LOGISIM_NET_93),
                        .pre(s_LOGISIM_NET_168));

   REGISTER_FLIP_FLOP_s6 #(.ActiveLevel(1),
                           .NrOfBits(32))
      REGISTER_FILE_32 (.Clock(LOGISIM_CLOCK_TREE_0[4]),
                        .ClockEnable(s_LOGISIM_NET_104),
                        .D(s_LOGISIM_BUS_136[31:0]),
                        .Q(s_LOGISIM_BUS_125[31:0]),
                        .Reset(s_LOGISIM_NET_34),
                        .Tick(LOGISIM_CLOCK_TREE_0[2]),
                        .cs(s_LOGISIM_NET_80),
                        .pre(s_LOGISIM_NET_167));

   Multiplexer_bus_32 #(.NrOfBits(32))
      MUX_2 (.Enable(1'b1),
             .MuxIn_0(s_LOGISIM_BUS_135[31:0]),
             .MuxIn_1(s_LOGISIM_BUS_56[31:0]),
             .MuxIn_10(s_LOGISIM_BUS_110[31:0]),
             .MuxIn_11(s_LOGISIM_BUS_124[31:0]),
             .MuxIn_12(s_LOGISIM_BUS_101[31:0]),
             .MuxIn_13(s_LOGISIM_BUS_18[31:0]),
             .MuxIn_14(s_LOGISIM_BUS_48[31:0]),
             .MuxIn_15(s_LOGISIM_BUS_108[31:0]),
             .MuxIn_16(s_LOGISIM_BUS_134[31:0]),
             .MuxIn_17(s_LOGISIM_BUS_57[31:0]),
             .MuxIn_18(s_LOGISIM_BUS_87[31:0]),
             .MuxIn_19(s_LOGISIM_BUS_85[31:0]),
             .MuxIn_2(s_LOGISIM_BUS_88[31:0]),
             .MuxIn_20(s_LOGISIM_BUS_100[31:0]),
             .MuxIn_21(s_LOGISIM_BUS_116[31:0]),
             .MuxIn_22(s_LOGISIM_BUS_132[31:0]),
             .MuxIn_23(s_LOGISIM_BUS_37[31:0]),
             .MuxIn_24(s_LOGISIM_BUS_67[31:0]),
             .MuxIn_25(s_LOGISIM_BUS_123[31:0]),
             .MuxIn_26(s_LOGISIM_BUS_66[31:0]),
             .MuxIn_27(s_LOGISIM_BUS_86[31:0]),
             .MuxIn_28(s_LOGISIM_BUS_102[31:0]),
             .MuxIn_29(s_LOGISIM_BUS_117[31:0]),
             .MuxIn_3(s_LOGISIM_BUS_76[31:0]),
             .MuxIn_30(s_LOGISIM_BUS_133[31:0]),
             .MuxIn_31(s_LOGISIM_BUS_109[31:0]),
             .MuxIn_4(s_LOGISIM_BUS_94[31:0]),
             .MuxIn_5(s_LOGISIM_BUS_111[31:0]),
             .MuxIn_6(s_LOGISIM_BUS_125[31:0]),
             .MuxIn_7(s_LOGISIM_BUS_36[31:0]),
             .MuxIn_8(s_LOGISIM_BUS_75[31:0]),
             .MuxIn_9(s_LOGISIM_BUS_122[31:0]),
             .MuxOut(s_LOGISIM_BUS_6[31:0]),
             .Sel(s_LOGISIM_BUS_26[4:0]));



endmodule
