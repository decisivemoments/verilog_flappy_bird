/******************************************************************************
 ** Logisim goes FPGA automatic generated Verilog code                       **
 **                                                                          **
 ** Component : signal_generator                                             **
 **                                                                          **
 ******************************************************************************/

`timescale 1ns/1ps
module signal_generator( F12,
                         F13,
                         F14,
                         F25,
                         F30,
                         LOGISIM_CLOCK_TREE_0,
                         OP2,
                         OP3,
                         OP4,
                         OP5,
                         OP6,
                         ALU_SRC,
                         AUIPC,
                         BEQ,
                         BLT,
                         BNE,
                         CSRRCI,
                         CSRRSI,
                         JAL,
                         JALR,
                         LBU,
                         MemToReg,
                         MemWrite,
                         RegWrite,
                         SRA,
                         S_Type,
                         ecall,
                         r1_used,
                         r2_used);

   /***************************************************************************
    ** Here the inputs are defined                                           **
    ***************************************************************************/
   input  F12;
   input  F13;
   input  F14;
   input  F25;
   input  F30;
   input[4:0]  LOGISIM_CLOCK_TREE_0;
   input  OP2;
   input  OP3;
   input  OP4;
   input  OP5;
   input  OP6;

   /***************************************************************************
    ** Here the outputs are defined                                          **
    ***************************************************************************/
   output ALU_SRC;
   output AUIPC;
   output BEQ;
   output BLT;
   output BNE;
   output CSRRCI;
   output CSRRSI;
   output JAL;
   output JALR;
   output LBU;
   output MemToReg;
   output MemWrite;
   output RegWrite;
   output SRA;
   output S_Type;
   output ecall;
   output r1_used;
   output r2_used;

   /***************************************************************************
    ** Here the internal wires are defined                                   **
    ***************************************************************************/
   wire s_LOGISIM_NET_0;
   wire s_LOGISIM_NET_1;
   wire s_LOGISIM_NET_10;
   wire s_LOGISIM_NET_100;
   wire s_LOGISIM_NET_101;
   wire s_LOGISIM_NET_102;
   wire s_LOGISIM_NET_103;
   wire s_LOGISIM_NET_104;
   wire s_LOGISIM_NET_105;
   wire s_LOGISIM_NET_106;
   wire s_LOGISIM_NET_107;
   wire s_LOGISIM_NET_108;
   wire s_LOGISIM_NET_109;
   wire s_LOGISIM_NET_11;
   wire s_LOGISIM_NET_110;
   wire s_LOGISIM_NET_111;
   wire s_LOGISIM_NET_112;
   wire s_LOGISIM_NET_113;
   wire s_LOGISIM_NET_114;
   wire s_LOGISIM_NET_115;
   wire s_LOGISIM_NET_116;
   wire s_LOGISIM_NET_117;
   wire s_LOGISIM_NET_118;
   wire s_LOGISIM_NET_119;
   wire s_LOGISIM_NET_12;
   wire s_LOGISIM_NET_120;
   wire s_LOGISIM_NET_121;
   wire s_LOGISIM_NET_122;
   wire s_LOGISIM_NET_123;
   wire s_LOGISIM_NET_124;
   wire s_LOGISIM_NET_125;
   wire s_LOGISIM_NET_126;
   wire s_LOGISIM_NET_127;
   wire s_LOGISIM_NET_128;
   wire s_LOGISIM_NET_129;
   wire s_LOGISIM_NET_13;
   wire s_LOGISIM_NET_130;
   wire s_LOGISIM_NET_131;
   wire s_LOGISIM_NET_132;
   wire s_LOGISIM_NET_133;
   wire s_LOGISIM_NET_134;
   wire s_LOGISIM_NET_135;
   wire s_LOGISIM_NET_136;
   wire s_LOGISIM_NET_137;
   wire s_LOGISIM_NET_138;
   wire s_LOGISIM_NET_139;
   wire s_LOGISIM_NET_14;
   wire s_LOGISIM_NET_140;
   wire s_LOGISIM_NET_141;
   wire s_LOGISIM_NET_142;
   wire s_LOGISIM_NET_143;
   wire s_LOGISIM_NET_144;
   wire s_LOGISIM_NET_145;
   wire s_LOGISIM_NET_146;
   wire s_LOGISIM_NET_147;
   wire s_LOGISIM_NET_148;
   wire s_LOGISIM_NET_149;
   wire s_LOGISIM_NET_15;
   wire s_LOGISIM_NET_150;
   wire s_LOGISIM_NET_151;
   wire s_LOGISIM_NET_152;
   wire s_LOGISIM_NET_153;
   wire s_LOGISIM_NET_154;
   wire s_LOGISIM_NET_155;
   wire s_LOGISIM_NET_156;
   wire s_LOGISIM_NET_157;
   wire s_LOGISIM_NET_158;
   wire s_LOGISIM_NET_159;
   wire s_LOGISIM_NET_16;
   wire s_LOGISIM_NET_160;
   wire s_LOGISIM_NET_161;
   wire s_LOGISIM_NET_162;
   wire s_LOGISIM_NET_163;
   wire s_LOGISIM_NET_164;
   wire s_LOGISIM_NET_165;
   wire s_LOGISIM_NET_166;
   wire s_LOGISIM_NET_167;
   wire s_LOGISIM_NET_168;
   wire s_LOGISIM_NET_169;
   wire s_LOGISIM_NET_17;
   wire s_LOGISIM_NET_170;
   wire s_LOGISIM_NET_171;
   wire s_LOGISIM_NET_172;
   wire s_LOGISIM_NET_173;
   wire s_LOGISIM_NET_174;
   wire s_LOGISIM_NET_175;
   wire s_LOGISIM_NET_176;
   wire s_LOGISIM_NET_177;
   wire s_LOGISIM_NET_178;
   wire s_LOGISIM_NET_179;
   wire s_LOGISIM_NET_18;
   wire s_LOGISIM_NET_180;
   wire s_LOGISIM_NET_181;
   wire s_LOGISIM_NET_182;
   wire s_LOGISIM_NET_183;
   wire s_LOGISIM_NET_184;
   wire s_LOGISIM_NET_185;
   wire s_LOGISIM_NET_186;
   wire s_LOGISIM_NET_187;
   wire s_LOGISIM_NET_188;
   wire s_LOGISIM_NET_189;
   wire s_LOGISIM_NET_19;
   wire s_LOGISIM_NET_190;
   wire s_LOGISIM_NET_191;
   wire s_LOGISIM_NET_192;
   wire s_LOGISIM_NET_193;
   wire s_LOGISIM_NET_194;
   wire s_LOGISIM_NET_195;
   wire s_LOGISIM_NET_196;
   wire s_LOGISIM_NET_197;
   wire s_LOGISIM_NET_198;
   wire s_LOGISIM_NET_199;
   wire s_LOGISIM_NET_2;
   wire s_LOGISIM_NET_20;
   wire s_LOGISIM_NET_200;
   wire s_LOGISIM_NET_201;
   wire s_LOGISIM_NET_202;
   wire s_LOGISIM_NET_203;
   wire s_LOGISIM_NET_204;
   wire s_LOGISIM_NET_205;
   wire s_LOGISIM_NET_206;
   wire s_LOGISIM_NET_207;
   wire s_LOGISIM_NET_208;
   wire s_LOGISIM_NET_209;
   wire s_LOGISIM_NET_21;
   wire s_LOGISIM_NET_210;
   wire s_LOGISIM_NET_211;
   wire s_LOGISIM_NET_212;
   wire s_LOGISIM_NET_213;
   wire s_LOGISIM_NET_214;
   wire s_LOGISIM_NET_215;
   wire s_LOGISIM_NET_216;
   wire s_LOGISIM_NET_217;
   wire s_LOGISIM_NET_218;
   wire s_LOGISIM_NET_219;
   wire s_LOGISIM_NET_22;
   wire s_LOGISIM_NET_220;
   wire s_LOGISIM_NET_221;
   wire s_LOGISIM_NET_222;
   wire s_LOGISIM_NET_223;
   wire s_LOGISIM_NET_224;
   wire s_LOGISIM_NET_225;
   wire s_LOGISIM_NET_226;
   wire s_LOGISIM_NET_227;
   wire s_LOGISIM_NET_228;
   wire s_LOGISIM_NET_229;
   wire s_LOGISIM_NET_23;
   wire s_LOGISIM_NET_230;
   wire s_LOGISIM_NET_231;
   wire s_LOGISIM_NET_232;
   wire s_LOGISIM_NET_233;
   wire s_LOGISIM_NET_234;
   wire s_LOGISIM_NET_235;
   wire s_LOGISIM_NET_236;
   wire s_LOGISIM_NET_237;
   wire s_LOGISIM_NET_238;
   wire s_LOGISIM_NET_239;
   wire s_LOGISIM_NET_24;
   wire s_LOGISIM_NET_240;
   wire s_LOGISIM_NET_241;
   wire s_LOGISIM_NET_242;
   wire s_LOGISIM_NET_243;
   wire s_LOGISIM_NET_244;
   wire s_LOGISIM_NET_245;
   wire s_LOGISIM_NET_246;
   wire s_LOGISIM_NET_247;
   wire s_LOGISIM_NET_248;
   wire s_LOGISIM_NET_249;
   wire s_LOGISIM_NET_25;
   wire s_LOGISIM_NET_250;
   wire s_LOGISIM_NET_251;
   wire s_LOGISIM_NET_252;
   wire s_LOGISIM_NET_253;
   wire s_LOGISIM_NET_254;
   wire s_LOGISIM_NET_255;
   wire s_LOGISIM_NET_256;
   wire s_LOGISIM_NET_257;
   wire s_LOGISIM_NET_258;
   wire s_LOGISIM_NET_259;
   wire s_LOGISIM_NET_26;
   wire s_LOGISIM_NET_260;
   wire s_LOGISIM_NET_261;
   wire s_LOGISIM_NET_262;
   wire s_LOGISIM_NET_263;
   wire s_LOGISIM_NET_264;
   wire s_LOGISIM_NET_265;
   wire s_LOGISIM_NET_266;
   wire s_LOGISIM_NET_267;
   wire s_LOGISIM_NET_268;
   wire s_LOGISIM_NET_269;
   wire s_LOGISIM_NET_27;
   wire s_LOGISIM_NET_270;
   wire s_LOGISIM_NET_271;
   wire s_LOGISIM_NET_272;
   wire s_LOGISIM_NET_273;
   wire s_LOGISIM_NET_274;
   wire s_LOGISIM_NET_275;
   wire s_LOGISIM_NET_276;
   wire s_LOGISIM_NET_277;
   wire s_LOGISIM_NET_278;
   wire s_LOGISIM_NET_279;
   wire s_LOGISIM_NET_28;
   wire s_LOGISIM_NET_280;
   wire s_LOGISIM_NET_281;
   wire s_LOGISIM_NET_282;
   wire s_LOGISIM_NET_283;
   wire s_LOGISIM_NET_284;
   wire s_LOGISIM_NET_285;
   wire s_LOGISIM_NET_286;
   wire s_LOGISIM_NET_287;
   wire s_LOGISIM_NET_288;
   wire s_LOGISIM_NET_289;
   wire s_LOGISIM_NET_29;
   wire s_LOGISIM_NET_290;
   wire s_LOGISIM_NET_291;
   wire s_LOGISIM_NET_292;
   wire s_LOGISIM_NET_293;
   wire s_LOGISIM_NET_294;
   wire s_LOGISIM_NET_295;
   wire s_LOGISIM_NET_296;
   wire s_LOGISIM_NET_297;
   wire s_LOGISIM_NET_298;
   wire s_LOGISIM_NET_299;
   wire s_LOGISIM_NET_3;
   wire s_LOGISIM_NET_30;
   wire s_LOGISIM_NET_300;
   wire s_LOGISIM_NET_301;
   wire s_LOGISIM_NET_302;
   wire s_LOGISIM_NET_303;
   wire s_LOGISIM_NET_304;
   wire s_LOGISIM_NET_305;
   wire s_LOGISIM_NET_306;
   wire s_LOGISIM_NET_307;
   wire s_LOGISIM_NET_308;
   wire s_LOGISIM_NET_309;
   wire s_LOGISIM_NET_31;
   wire s_LOGISIM_NET_310;
   wire s_LOGISIM_NET_311;
   wire s_LOGISIM_NET_312;
   wire s_LOGISIM_NET_313;
   wire s_LOGISIM_NET_314;
   wire s_LOGISIM_NET_315;
   wire s_LOGISIM_NET_316;
   wire s_LOGISIM_NET_317;
   wire s_LOGISIM_NET_318;
   wire s_LOGISIM_NET_319;
   wire s_LOGISIM_NET_32;
   wire s_LOGISIM_NET_320;
   wire s_LOGISIM_NET_321;
   wire s_LOGISIM_NET_322;
   wire s_LOGISIM_NET_323;
   wire s_LOGISIM_NET_324;
   wire s_LOGISIM_NET_325;
   wire s_LOGISIM_NET_326;
   wire s_LOGISIM_NET_327;
   wire s_LOGISIM_NET_328;
   wire s_LOGISIM_NET_329;
   wire s_LOGISIM_NET_33;
   wire s_LOGISIM_NET_330;
   wire s_LOGISIM_NET_331;
   wire s_LOGISIM_NET_332;
   wire s_LOGISIM_NET_333;
   wire s_LOGISIM_NET_334;
   wire s_LOGISIM_NET_335;
   wire s_LOGISIM_NET_336;
   wire s_LOGISIM_NET_337;
   wire s_LOGISIM_NET_338;
   wire s_LOGISIM_NET_339;
   wire s_LOGISIM_NET_34;
   wire s_LOGISIM_NET_340;
   wire s_LOGISIM_NET_341;
   wire s_LOGISIM_NET_342;
   wire s_LOGISIM_NET_343;
   wire s_LOGISIM_NET_344;
   wire s_LOGISIM_NET_345;
   wire s_LOGISIM_NET_346;
   wire s_LOGISIM_NET_347;
   wire s_LOGISIM_NET_348;
   wire s_LOGISIM_NET_349;
   wire s_LOGISIM_NET_35;
   wire s_LOGISIM_NET_350;
   wire s_LOGISIM_NET_351;
   wire s_LOGISIM_NET_352;
   wire s_LOGISIM_NET_353;
   wire s_LOGISIM_NET_354;
   wire s_LOGISIM_NET_355;
   wire s_LOGISIM_NET_356;
   wire s_LOGISIM_NET_357;
   wire s_LOGISIM_NET_358;
   wire s_LOGISIM_NET_359;
   wire s_LOGISIM_NET_36;
   wire s_LOGISIM_NET_360;
   wire s_LOGISIM_NET_361;
   wire s_LOGISIM_NET_362;
   wire s_LOGISIM_NET_363;
   wire s_LOGISIM_NET_364;
   wire s_LOGISIM_NET_365;
   wire s_LOGISIM_NET_366;
   wire s_LOGISIM_NET_367;
   wire s_LOGISIM_NET_368;
   wire s_LOGISIM_NET_369;
   wire s_LOGISIM_NET_37;
   wire s_LOGISIM_NET_370;
   wire s_LOGISIM_NET_371;
   wire s_LOGISIM_NET_372;
   wire s_LOGISIM_NET_373;
   wire s_LOGISIM_NET_374;
   wire s_LOGISIM_NET_375;
   wire s_LOGISIM_NET_376;
   wire s_LOGISIM_NET_377;
   wire s_LOGISIM_NET_378;
   wire s_LOGISIM_NET_379;
   wire s_LOGISIM_NET_38;
   wire s_LOGISIM_NET_380;
   wire s_LOGISIM_NET_381;
   wire s_LOGISIM_NET_382;
   wire s_LOGISIM_NET_383;
   wire s_LOGISIM_NET_384;
   wire s_LOGISIM_NET_385;
   wire s_LOGISIM_NET_386;
   wire s_LOGISIM_NET_387;
   wire s_LOGISIM_NET_388;
   wire s_LOGISIM_NET_389;
   wire s_LOGISIM_NET_39;
   wire s_LOGISIM_NET_390;
   wire s_LOGISIM_NET_391;
   wire s_LOGISIM_NET_392;
   wire s_LOGISIM_NET_393;
   wire s_LOGISIM_NET_394;
   wire s_LOGISIM_NET_395;
   wire s_LOGISIM_NET_396;
   wire s_LOGISIM_NET_397;
   wire s_LOGISIM_NET_398;
   wire s_LOGISIM_NET_399;
   wire s_LOGISIM_NET_4;
   wire s_LOGISIM_NET_40;
   wire s_LOGISIM_NET_400;
   wire s_LOGISIM_NET_401;
   wire s_LOGISIM_NET_402;
   wire s_LOGISIM_NET_403;
   wire s_LOGISIM_NET_41;
   wire s_LOGISIM_NET_42;
   wire s_LOGISIM_NET_43;
   wire s_LOGISIM_NET_44;
   wire s_LOGISIM_NET_45;
   wire s_LOGISIM_NET_46;
   wire s_LOGISIM_NET_47;
   wire s_LOGISIM_NET_48;
   wire s_LOGISIM_NET_49;
   wire s_LOGISIM_NET_5;
   wire s_LOGISIM_NET_50;
   wire s_LOGISIM_NET_51;
   wire s_LOGISIM_NET_52;
   wire s_LOGISIM_NET_53;
   wire s_LOGISIM_NET_54;
   wire s_LOGISIM_NET_55;
   wire s_LOGISIM_NET_56;
   wire s_LOGISIM_NET_57;
   wire s_LOGISIM_NET_58;
   wire s_LOGISIM_NET_59;
   wire s_LOGISIM_NET_6;
   wire s_LOGISIM_NET_60;
   wire s_LOGISIM_NET_61;
   wire s_LOGISIM_NET_62;
   wire s_LOGISIM_NET_63;
   wire s_LOGISIM_NET_64;
   wire s_LOGISIM_NET_65;
   wire s_LOGISIM_NET_66;
   wire s_LOGISIM_NET_67;
   wire s_LOGISIM_NET_68;
   wire s_LOGISIM_NET_69;
   wire s_LOGISIM_NET_7;
   wire s_LOGISIM_NET_70;
   wire s_LOGISIM_NET_71;
   wire s_LOGISIM_NET_72;
   wire s_LOGISIM_NET_73;
   wire s_LOGISIM_NET_74;
   wire s_LOGISIM_NET_75;
   wire s_LOGISIM_NET_76;
   wire s_LOGISIM_NET_77;
   wire s_LOGISIM_NET_78;
   wire s_LOGISIM_NET_79;
   wire s_LOGISIM_NET_8;
   wire s_LOGISIM_NET_80;
   wire s_LOGISIM_NET_81;
   wire s_LOGISIM_NET_82;
   wire s_LOGISIM_NET_83;
   wire s_LOGISIM_NET_84;
   wire s_LOGISIM_NET_85;
   wire s_LOGISIM_NET_86;
   wire s_LOGISIM_NET_87;
   wire s_LOGISIM_NET_88;
   wire s_LOGISIM_NET_89;
   wire s_LOGISIM_NET_9;
   wire s_LOGISIM_NET_90;
   wire s_LOGISIM_NET_91;
   wire s_LOGISIM_NET_92;
   wire s_LOGISIM_NET_93;
   wire s_LOGISIM_NET_94;
   wire s_LOGISIM_NET_95;
   wire s_LOGISIM_NET_96;
   wire s_LOGISIM_NET_97;
   wire s_LOGISIM_NET_98;
   wire s_LOGISIM_NET_99;


   /***************************************************************************
    ** Here all input connections are defined                                **
    ***************************************************************************/
   assign s_LOGISIM_NET_18                   = F30;
   assign s_LOGISIM_NET_7                    = F13;
   assign s_LOGISIM_NET_5                    = F14;
   assign s_LOGISIM_NET_22                   = OP3;
   assign s_LOGISIM_NET_10                   = F25;
   assign s_LOGISIM_NET_35                   = F12;
   assign s_LOGISIM_NET_31                   = OP6;
   assign s_LOGISIM_NET_9                    = OP4;
   assign s_LOGISIM_NET_14                   = OP2;
   assign s_LOGISIM_NET_32                   = OP5;

   /***************************************************************************
    ** Here all output connections are defined                               **
    ***************************************************************************/
   assign RegWrite                           = s_LOGISIM_NET_389;
   assign CSRRCI                             = s_LOGISIM_NET_394;
   assign ALU_SRC                            = s_LOGISIM_NET_359;
   assign JAL                                = s_LOGISIM_NET_381;
   assign CSRRSI                             = s_LOGISIM_NET_373;
   assign SRA                                = s_LOGISIM_NET_399;
   assign S_Type                             = s_LOGISIM_NET_392;
   assign BLT                                = s_LOGISIM_NET_369;
   assign r2_used                            = s_LOGISIM_NET_383;
   assign LBU                                = s_LOGISIM_NET_26;
   assign r1_used                            = s_LOGISIM_NET_372;
   assign BEQ                                = s_LOGISIM_NET_284;
   assign MemToReg                           = s_LOGISIM_NET_377;
   assign AUIPC                              = s_LOGISIM_NET_401;
   assign MemWrite                           = s_LOGISIM_NET_386;
   assign JALR                               = s_LOGISIM_NET_268;
   assign BNE                                = s_LOGISIM_NET_2;
   assign ecall                              = s_LOGISIM_NET_184;

   /***************************************************************************
    ** Here all normal components are defined                                **
    ***************************************************************************/
   NOT_GATE      GATE_1 (.Input_1(s_LOGISIM_NET_7),
                         .Result(s_LOGISIM_NET_54));

   AND_GATE_8_INPUTS #(.BubblesMask(0))
      GATE_2 (.Input_1(s_LOGISIM_NET_14),
              .Input_2(s_LOGISIM_NET_279),
              .Input_3(s_LOGISIM_NET_93),
              .Input_4(s_LOGISIM_NET_32),
              .Input_5(s_LOGISIM_NET_31),
              .Input_6(s_LOGISIM_NET_102),
              .Input_7(s_LOGISIM_NET_320),
              .Input_8(s_LOGISIM_NET_114),
              .Result(s_LOGISIM_NET_268));

   NOT_GATE      GATE_3 (.Input_1(s_LOGISIM_NET_14),
                         .Result(s_LOGISIM_NET_92));

   NOT_GATE      GATE_4 (.Input_1(s_LOGISIM_NET_14),
                         .Result(s_LOGISIM_NET_110));

   AND_GATE_10_INPUTS #(.BubblesMask(0))
      GATE_5 (.Input_1(s_LOGISIM_NET_156),
              .Input_10(s_LOGISIM_NET_18),
              .Input_2(s_LOGISIM_NET_339),
              .Input_3(s_LOGISIM_NET_9),
              .Input_4(s_LOGISIM_NET_32),
              .Input_5(s_LOGISIM_NET_300),
              .Input_6(s_LOGISIM_NET_35),
              .Input_7(s_LOGISIM_NET_240),
              .Input_8(s_LOGISIM_NET_5),
              .Input_9(s_LOGISIM_NET_244),
              .Result(s_LOGISIM_NET_399));

   AND_GATE_5_INPUTS #(.BubblesMask(0))
      GATE_6 (.Input_1(s_LOGISIM_NET_40),
              .Input_2(s_LOGISIM_NET_325),
              .Input_3(s_LOGISIM_NET_9),
              .Input_4(s_LOGISIM_NET_86),
              .Input_5(s_LOGISIM_NET_14),
              .Result(s_LOGISIM_NET_361));

   NOT_GATE      GATE_7 (.Input_1(s_LOGISIM_NET_35),
                         .Result(s_LOGISIM_NET_171));

   NOT_GATE      GATE_8 (.Input_1(s_LOGISIM_NET_14),
                         .Result(s_LOGISIM_NET_76));

   AND_GATE_7_INPUTS #(.BubblesMask(0))
      GATE_9 (.Input_1(s_LOGISIM_NET_192),
              .Input_2(s_LOGISIM_NET_6),
              .Input_3(s_LOGISIM_NET_124),
              .Input_4(s_LOGISIM_NET_32),
              .Input_5(s_LOGISIM_NET_31),
              .Input_6(s_LOGISIM_NET_351),
              .Input_7(s_LOGISIM_NET_70),
              .Result(s_LOGISIM_NET_158));

   NOT_GATE      GATE_10 (.Input_1(s_LOGISIM_NET_31),
                          .Result(s_LOGISIM_NET_328));

   NOT_GATE      GATE_11 (.Input_1(s_LOGISIM_NET_14),
                          .Result(s_LOGISIM_NET_224));

   NOT_GATE      GATE_12 (.Input_1(s_LOGISIM_NET_35),
                          .Result(s_LOGISIM_NET_338));

   NOT_GATE      GATE_13 (.Input_1(s_LOGISIM_NET_14),
                          .Result(s_LOGISIM_NET_21));

   NOT_GATE      GATE_14 (.Input_1(s_LOGISIM_NET_7),
                          .Result(s_LOGISIM_NET_185));

   NOT_GATE      GATE_15 (.Input_1(s_LOGISIM_NET_22),
                          .Result(s_LOGISIM_NET_122));

   NOT_GATE      GATE_16 (.Input_1(s_LOGISIM_NET_35),
                          .Result(s_LOGISIM_NET_62));

   AND_GATE_8_INPUTS #(.BubblesMask(0))
      GATE_17 (.Input_1(s_LOGISIM_NET_5),
               .Input_2(s_LOGISIM_NET_172),
               .Input_3(s_LOGISIM_NET_312),
               .Input_4(s_LOGISIM_NET_327),
               .Input_5(s_LOGISIM_NET_262),
               .Input_6(s_LOGISIM_NET_319),
               .Input_7(s_LOGISIM_NET_169),
               .Input_8(s_LOGISIM_NET_224),
               .Result(s_LOGISIM_NET_41));

   NOT_GATE      GATE_18 (.Input_1(s_LOGISIM_NET_35),
                          .Result(s_LOGISIM_NET_89));

   AND_GATE_7_INPUTS #(.BubblesMask(0))
      GATE_19 (.Input_1(s_LOGISIM_NET_337),
               .Input_2(s_LOGISIM_NET_219),
               .Input_3(s_LOGISIM_NET_340),
               .Input_4(s_LOGISIM_NET_285),
               .Input_5(s_LOGISIM_NET_134),
               .Input_6(s_LOGISIM_NET_273),
               .Input_7(s_LOGISIM_NET_5),
               .Result(s_LOGISIM_NET_164));

   NOT_GATE      GATE_20 (.Input_1(s_LOGISIM_NET_14),
                          .Result(s_LOGISIM_NET_23));

   NOT_GATE      GATE_21 (.Input_1(s_LOGISIM_NET_9),
                          .Result(s_LOGISIM_NET_334));

   NOT_GATE      GATE_22 (.Input_1(s_LOGISIM_NET_31),
                          .Result(s_LOGISIM_NET_384));

   NOT_GATE      GATE_23 (.Input_1(s_LOGISIM_NET_7),
                          .Result(s_LOGISIM_NET_203));

   NOT_GATE      GATE_24 (.Input_1(s_LOGISIM_NET_22),
                          .Result(s_LOGISIM_NET_84));

   NOT_GATE      GATE_25 (.Input_1(s_LOGISIM_NET_31),
                          .Result(s_LOGISIM_NET_403));

   NOT_GATE      GATE_26 (.Input_1(s_LOGISIM_NET_32),
                          .Result(s_LOGISIM_NET_402));

   NOT_GATE      GATE_27 (.Input_1(s_LOGISIM_NET_22),
                          .Result(s_LOGISIM_NET_219));

   NOT_GATE      GATE_28 (.Input_1(s_LOGISIM_NET_22),
                          .Result(s_LOGISIM_NET_135));

   OR_GATE_7_INPUTS #(.BubblesMask(0))
      GATE_29 (.Input_1(s_LOGISIM_NET_188),
               .Input_2(s_LOGISIM_NET_290),
               .Input_3(s_LOGISIM_NET_104),
               .Input_4(s_LOGISIM_NET_333),
               .Input_5(s_LOGISIM_NET_3),
               .Input_6(s_LOGISIM_NET_207),
               .Input_7(s_LOGISIM_NET_87),
               .Result(s_LOGISIM_NET_359));

   NOT_GATE      GATE_30 (.Input_1(s_LOGISIM_NET_22),
                          .Result(s_LOGISIM_NET_37));

   NOT_GATE      GATE_31 (.Input_1(s_LOGISIM_NET_10),
                          .Result(s_LOGISIM_NET_1));

   NOT_GATE      GATE_32 (.Input_1(s_LOGISIM_NET_14),
                          .Result(s_LOGISIM_NET_258));

   NOT_GATE      GATE_33 (.Input_1(s_LOGISIM_NET_14),
                          .Result(s_LOGISIM_NET_45));

   NOT_GATE      GATE_34 (.Input_1(s_LOGISIM_NET_9),
                          .Result(s_LOGISIM_NET_296));

   AND_GATE_8_INPUTS #(.BubblesMask(0))
      GATE_35 (.Input_1(s_LOGISIM_NET_162),
               .Input_2(s_LOGISIM_NET_7),
               .Input_3(s_LOGISIM_NET_83),
               .Input_4(s_LOGISIM_NET_115),
               .Input_5(s_LOGISIM_NET_357),
               .Input_6(s_LOGISIM_NET_9),
               .Input_7(s_LOGISIM_NET_311),
               .Input_8(s_LOGISIM_NET_99),
               .Result(s_LOGISIM_NET_398));

   NOT_GATE      GATE_36 (.Input_1(s_LOGISIM_NET_31),
                          .Result(s_LOGISIM_NET_378));

   NOT_GATE      GATE_37 (.Input_1(s_LOGISIM_NET_32),
                          .Result(s_LOGISIM_NET_229));

   NOT_GATE      GATE_38 (.Input_1(s_LOGISIM_NET_35),
                          .Result(s_LOGISIM_NET_29));

   NOT_GATE      GATE_39 (.Input_1(s_LOGISIM_NET_9),
                          .Result(s_LOGISIM_NET_289));

   NOT_GATE      GATE_40 (.Input_1(s_LOGISIM_NET_5),
                          .Result(s_LOGISIM_NET_59));

   NOT_GATE      GATE_41 (.Input_1(s_LOGISIM_NET_9),
                          .Result(s_LOGISIM_NET_319));

   NOT_GATE      GATE_42 (.Input_1(s_LOGISIM_NET_7),
                          .Result(s_LOGISIM_NET_106));

   NOT_GATE      GATE_43 (.Input_1(s_LOGISIM_NET_31),
                          .Result(s_LOGISIM_NET_395));

   NOT_GATE      GATE_44 (.Input_1(s_LOGISIM_NET_18),
                          .Result(s_LOGISIM_NET_209));

   NOT_GATE      GATE_45 (.Input_1(s_LOGISIM_NET_7),
                          .Result(s_LOGISIM_NET_68));

   NOT_GATE      GATE_46 (.Input_1(s_LOGISIM_NET_9),
                          .Result(s_LOGISIM_NET_121));

   AND_GATE_8_INPUTS #(.BubblesMask(0))
      GATE_47 (.Input_1(s_LOGISIM_NET_144),
               .Input_2(s_LOGISIM_NET_36),
               .Input_3(s_LOGISIM_NET_182),
               .Input_4(s_LOGISIM_NET_31),
               .Input_5(s_LOGISIM_NET_32),
               .Input_6(s_LOGISIM_NET_362),
               .Input_7(s_LOGISIM_NET_123),
               .Input_8(s_LOGISIM_NET_14),
               .Result(s_LOGISIM_NET_356));

   AND_GATE_10_INPUTS #(.BubblesMask(0))
      GATE_48 (.Input_1(s_LOGISIM_NET_237),
               .Input_10(s_LOGISIM_NET_77),
               .Input_2(s_LOGISIM_NET_12),
               .Input_3(s_LOGISIM_NET_5),
               .Input_4(s_LOGISIM_NET_28),
               .Input_5(s_LOGISIM_NET_35),
               .Input_6(s_LOGISIM_NET_371),
               .Input_7(s_LOGISIM_NET_305),
               .Input_8(s_LOGISIM_NET_9),
               .Input_9(s_LOGISIM_NET_306),
               .Result(s_LOGISIM_NET_69));

   NOT_GATE      GATE_49 (.Input_1(s_LOGISIM_NET_9),
                          .Result(s_LOGISIM_NET_343));

   AND_GATE_7_INPUTS #(.BubblesMask(0))
      GATE_50 (.Input_1(s_LOGISIM_NET_303),
               .Input_2(s_LOGISIM_NET_145),
               .Input_3(s_LOGISIM_NET_334),
               .Input_4(s_LOGISIM_NET_32),
               .Input_5(s_LOGISIM_NET_31),
               .Input_6(s_LOGISIM_NET_201),
               .Input_7(s_LOGISIM_NET_353),
               .Result(s_LOGISIM_NET_177));

   NOT_GATE      GATE_51 (.Input_1(s_LOGISIM_NET_32),
                          .Result(s_LOGISIM_NET_325));

   AND_GATE_9_INPUTS #(.BubblesMask(0))
      GATE_52 (.Input_1(s_LOGISIM_NET_215),
               .Input_2(s_LOGISIM_NET_74),
               .Input_3(s_LOGISIM_NET_9),
               .Input_4(s_LOGISIM_NET_32),
               .Input_5(s_LOGISIM_NET_238),
               .Input_6(s_LOGISIM_NET_62),
               .Input_7(s_LOGISIM_NET_181),
               .Input_8(s_LOGISIM_NET_376),
               .Input_9(s_LOGISIM_NET_80),
               .Result(s_LOGISIM_NET_127));

   NOT_GATE      GATE_53 (.Input_1(s_LOGISIM_NET_31),
                          .Result(s_LOGISIM_NET_246));

   NOT_GATE      GATE_54 (.Input_1(s_LOGISIM_NET_31),
                          .Result(s_LOGISIM_NET_302));

   NOT_GATE      GATE_55 (.Input_1(s_LOGISIM_NET_9),
                          .Result(s_LOGISIM_NET_8));

   NOT_GATE      GATE_56 (.Input_1(s_LOGISIM_NET_31),
                          .Result(s_LOGISIM_NET_238));

   NOT_GATE      GATE_57 (.Input_1(s_LOGISIM_NET_31),
                          .Result(s_LOGISIM_NET_226));

   NOT_GATE      GATE_58 (.Input_1(s_LOGISIM_NET_14),
                          .Result(s_LOGISIM_NET_282));

   NOT_GATE      GATE_59 (.Input_1(s_LOGISIM_NET_35),
                          .Result(s_LOGISIM_NET_264));

   AND_GATE_10_INPUTS #(.BubblesMask(0))
      GATE_60 (.Input_1(s_LOGISIM_NET_150),
               .Input_10(s_LOGISIM_NET_332),
               .Input_2(s_LOGISIM_NET_10),
               .Input_3(s_LOGISIM_NET_254),
               .Input_4(s_LOGISIM_NET_50),
               .Input_5(s_LOGISIM_NET_89),
               .Input_6(s_LOGISIM_NET_328),
               .Input_7(s_LOGISIM_NET_32),
               .Input_8(s_LOGISIM_NET_9),
               .Input_9(s_LOGISIM_NET_190),
               .Result(s_LOGISIM_NET_34));

   NOT_GATE      GATE_61 (.Input_1(s_LOGISIM_NET_14),
                          .Result(s_LOGISIM_NET_337));

   AND_GATE_7_INPUTS #(.BubblesMask(0))
      GATE_62 (.Input_1(s_LOGISIM_NET_101),
               .Input_2(s_LOGISIM_NET_314),
               .Input_3(s_LOGISIM_NET_13),
               .Input_4(s_LOGISIM_NET_350),
               .Input_5(s_LOGISIM_NET_29),
               .Input_6(s_LOGISIM_NET_341),
               .Input_7(s_LOGISIM_NET_5),
               .Result(s_LOGISIM_NET_188));

   NOT_GATE      GATE_63 (.Input_1(s_LOGISIM_NET_18),
                          .Result(s_LOGISIM_NET_222));

   NOT_GATE      GATE_64 (.Input_1(s_LOGISIM_NET_18),
                          .Result(s_LOGISIM_NET_278));

   NOT_GATE      GATE_65 (.Input_1(s_LOGISIM_NET_31),
                          .Result(s_LOGISIM_NET_307));

   NOT_GATE      GATE_66 (.Input_1(s_LOGISIM_NET_31),
                          .Result(s_LOGISIM_NET_299));

   AND_GATE_10_INPUTS #(.BubblesMask(0))
      GATE_67 (.Input_1(s_LOGISIM_NET_21),
               .Input_10(s_LOGISIM_NET_140),
               .Input_2(s_LOGISIM_NET_175),
               .Input_3(s_LOGISIM_NET_9),
               .Input_4(s_LOGISIM_NET_32),
               .Input_5(s_LOGISIM_NET_31),
               .Input_6(s_LOGISIM_NET_400),
               .Input_7(s_LOGISIM_NET_364),
               .Input_8(s_LOGISIM_NET_56),
               .Input_9(s_LOGISIM_NET_277),
               .Result(s_LOGISIM_NET_184));

   AND_GATE_8_INPUTS #(.BubblesMask(0))
      GATE_68 (.Input_1(s_LOGISIM_NET_14),
               .Input_2(s_LOGISIM_NET_179),
               .Input_3(s_LOGISIM_NET_289),
               .Input_4(s_LOGISIM_NET_32),
               .Input_5(s_LOGISIM_NET_31),
               .Input_6(s_LOGISIM_NET_292),
               .Input_7(s_LOGISIM_NET_108),
               .Input_8(s_LOGISIM_NET_51),
               .Result(s_LOGISIM_NET_87));

   NOT_GATE      GATE_69 (.Input_1(s_LOGISIM_NET_31),
                          .Result(s_LOGISIM_NET_73));

   NOT_GATE      GATE_70 (.Input_1(s_LOGISIM_NET_31),
                          .Result(s_LOGISIM_NET_147));

   NOT_GATE      GATE_71 (.Input_1(s_LOGISIM_NET_14),
                          .Result(s_LOGISIM_NET_308));

   NOT_GATE      GATE_72 (.Input_1(s_LOGISIM_NET_14),
                          .Result(s_LOGISIM_NET_130));

   NOT_GATE      GATE_73 (.Input_1(s_LOGISIM_NET_32),
                          .Result(s_LOGISIM_NET_396));

   NOT_GATE      GATE_74 (.Input_1(s_LOGISIM_NET_5),
                          .Result(s_LOGISIM_NET_78));

   NOT_GATE      GATE_75 (.Input_1(s_LOGISIM_NET_35),
                          .Result(s_LOGISIM_NET_223));

   NOT_GATE      GATE_76 (.Input_1(s_LOGISIM_NET_7),
                          .Result(s_LOGISIM_NET_28));

   NOT_GATE      GATE_77 (.Input_1(s_LOGISIM_NET_22),
                          .Result(s_LOGISIM_NET_24));

   NOT_GATE      GATE_78 (.Input_1(s_LOGISIM_NET_5),
                          .Result(s_LOGISIM_NET_376));

   AND_GATE_10_INPUTS #(.BubblesMask(0))
      GATE_79 (.Input_1(s_LOGISIM_NET_278),
               .Input_10(s_LOGISIM_NET_143),
               .Input_2(s_LOGISIM_NET_95),
               .Input_3(s_LOGISIM_NET_5),
               .Input_4(s_LOGISIM_NET_7),
               .Input_5(s_LOGISIM_NET_360),
               .Input_6(s_LOGISIM_NET_291),
               .Input_7(s_LOGISIM_NET_32),
               .Input_8(s_LOGISIM_NET_9),
               .Input_9(s_LOGISIM_NET_336),
               .Result(s_LOGISIM_NET_91));

   NOT_GATE      GATE_80 (.Input_1(s_LOGISIM_NET_9),
                          .Result(s_LOGISIM_NET_142));

   NOT_GATE      GATE_81 (.Input_1(s_LOGISIM_NET_31),
                          .Result(s_LOGISIM_NET_371));

   NOT_GATE      GATE_82 (.Input_1(s_LOGISIM_NET_31),
                          .Result(s_LOGISIM_NET_199));

   NOT_GATE      GATE_83 (.Input_1(s_LOGISIM_NET_14),
                          .Result(s_LOGISIM_NET_216));

   NOT_GATE      GATE_84 (.Input_1(s_LOGISIM_NET_22),
                          .Result(s_LOGISIM_NET_86));

   NOT_GATE      GATE_85 (.Input_1(s_LOGISIM_NET_5),
                          .Result(s_LOGISIM_NET_144));

   NOT_GATE      GATE_86 (.Input_1(s_LOGISIM_NET_5),
                          .Result(s_LOGISIM_NET_212));

   NOT_GATE      GATE_87 (.Input_1(s_LOGISIM_NET_22),
                          .Result(s_LOGISIM_NET_248));

   NOT_GATE      GATE_88 (.Input_1(s_LOGISIM_NET_31),
                          .Result(s_LOGISIM_NET_397));

   NOT_GATE      GATE_89 (.Input_1(s_LOGISIM_NET_14),
                          .Result(s_LOGISIM_NET_25));

   AND_GATE_8_INPUTS #(.BubblesMask(0))
      GATE_90 (.Input_1(s_LOGISIM_NET_5),
               .Input_2(s_LOGISIM_NET_7),
               .Input_3(s_LOGISIM_NET_35),
               .Input_4(s_LOGISIM_NET_355),
               .Input_5(s_LOGISIM_NET_65),
               .Input_6(s_LOGISIM_NET_9),
               .Input_7(s_LOGISIM_NET_71),
               .Input_8(s_LOGISIM_NET_195),
               .Result(s_LOGISIM_NET_17));

   NOT_GATE      GATE_91 (.Input_1(s_LOGISIM_NET_22),
                          .Result(s_LOGISIM_NET_169));

   NOT_GATE      GATE_92 (.Input_1(s_LOGISIM_NET_22),
                          .Result(s_LOGISIM_NET_367));

   NOT_GATE      GATE_93 (.Input_1(s_LOGISIM_NET_32),
                          .Result(s_LOGISIM_NET_193));

   NOT_GATE      GATE_94 (.Input_1(s_LOGISIM_NET_7),
                          .Result(s_LOGISIM_NET_233));

   NOT_GATE      GATE_95 (.Input_1(s_LOGISIM_NET_32),
                          .Result(s_LOGISIM_NET_340));

   NOT_GATE      GATE_96 (.Input_1(s_LOGISIM_NET_14),
                          .Result(s_LOGISIM_NET_370));

   NOT_GATE      GATE_97 (.Input_1(s_LOGISIM_NET_10),
                          .Result(s_LOGISIM_NET_382));

   NOT_GATE      GATE_98 (.Input_1(s_LOGISIM_NET_7),
                          .Result(s_LOGISIM_NET_231));

   NOT_GATE      GATE_99 (.Input_1(s_LOGISIM_NET_7),
                          .Result(s_LOGISIM_NET_243));

   NOT_GATE      GATE_100 (.Input_1(s_LOGISIM_NET_10),
                           .Result(s_LOGISIM_NET_80));

   NOT_GATE      GATE_101 (.Input_1(s_LOGISIM_NET_22),
                           .Result(s_LOGISIM_NET_280));

   NOT_GATE      GATE_102 (.Input_1(s_LOGISIM_NET_22),
                           .Result(s_LOGISIM_NET_71));

   NOT_GATE      GATE_103 (.Input_1(s_LOGISIM_NET_9),
                           .Result(s_LOGISIM_NET_194));

   NOT_GATE      GATE_104 (.Input_1(s_LOGISIM_NET_10),
                           .Result(s_LOGISIM_NET_345));

   NOT_GATE      GATE_105 (.Input_1(s_LOGISIM_NET_7),
                           .Result(s_LOGISIM_NET_160));

   NOT_GATE      GATE_106 (.Input_1(s_LOGISIM_NET_5),
                           .Result(s_LOGISIM_NET_120));

   NOT_GATE      GATE_107 (.Input_1(s_LOGISIM_NET_10),
                           .Result(s_LOGISIM_NET_380));

   NOT_GATE      GATE_108 (.Input_1(s_LOGISIM_NET_22),
                           .Result(s_LOGISIM_NET_60));

   NOT_GATE      GATE_109 (.Input_1(s_LOGISIM_NET_18),
                           .Result(s_LOGISIM_NET_189));

   NOT_GATE      GATE_110 (.Input_1(s_LOGISIM_NET_22),
                           .Result(s_LOGISIM_NET_176));

   NOT_GATE      GATE_111 (.Input_1(s_LOGISIM_NET_31),
                           .Result(s_LOGISIM_NET_98));

   NOT_GATE      GATE_112 (.Input_1(s_LOGISIM_NET_22),
                           .Result(s_LOGISIM_NET_4));

   NOT_GATE      GATE_113 (.Input_1(s_LOGISIM_NET_31),
                           .Result(s_LOGISIM_NET_250));

   NOT_GATE      GATE_114 (.Input_1(s_LOGISIM_NET_22),
                           .Result(s_LOGISIM_NET_159));

   NOT_GATE      GATE_115 (.Input_1(s_LOGISIM_NET_22),
                           .Result(s_LOGISIM_NET_145));

   AND_GATE_8_INPUTS #(.BubblesMask(0))
      GATE_116 (.Input_1(s_LOGISIM_NET_130),
                .Input_2(s_LOGISIM_NET_297),
                .Input_3(s_LOGISIM_NET_121),
                .Input_4(s_LOGISIM_NET_32),
                .Input_5(s_LOGISIM_NET_31),
                .Input_6(s_LOGISIM_NET_132),
                .Input_7(s_LOGISIM_NET_330),
                .Input_8(s_LOGISIM_NET_148),
                .Result(s_LOGISIM_NET_284));

   NOT_GATE      GATE_117 (.Input_1(s_LOGISIM_NET_35),
                           .Result(s_LOGISIM_NET_344));

   NOT_GATE      GATE_118 (.Input_1(s_LOGISIM_NET_5),
                           .Result(s_LOGISIM_NET_118));

   NOT_GATE      GATE_119 (.Input_1(s_LOGISIM_NET_32),
                           .Result(s_LOGISIM_NET_305));

   NOT_GATE      GATE_120 (.Input_1(s_LOGISIM_NET_22),
                           .Result(s_LOGISIM_NET_16));

   AND_GATE_7_INPUTS #(.BubblesMask(0))
      GATE_121 (.Input_1(s_LOGISIM_NET_298),
                .Input_2(s_LOGISIM_NET_161),
                .Input_3(s_LOGISIM_NET_8),
                .Input_4(s_LOGISIM_NET_395),
                .Input_5(s_LOGISIM_NET_264),
                .Input_6(s_LOGISIM_NET_7),
                .Input_7(s_LOGISIM_NET_212),
                .Result(s_LOGISIM_NET_323));

   NOT_GATE      GATE_122 (.Input_1(s_LOGISIM_NET_22),
                           .Result(s_LOGISIM_NET_288));

   NOT_GATE      GATE_123 (.Input_1(s_LOGISIM_NET_7),
                           .Result(s_LOGISIM_NET_214));

   NOT_GATE      GATE_124 (.Input_1(s_LOGISIM_NET_32),
                           .Result(s_LOGISIM_NET_163));

   NOT_GATE      GATE_125 (.Input_1(s_LOGISIM_NET_9),
                           .Result(s_LOGISIM_NET_274));

   NOT_GATE      GATE_126 (.Input_1(s_LOGISIM_NET_32),
                           .Result(s_LOGISIM_NET_109));

   NOT_GATE      GATE_127 (.Input_1(s_LOGISIM_NET_14),
                           .Result(s_LOGISIM_NET_61));

   NOT_GATE      GATE_128 (.Input_1(s_LOGISIM_NET_5),
                           .Result(s_LOGISIM_NET_51));

   NOT_GATE      GATE_129 (.Input_1(s_LOGISIM_NET_22),
                           .Result(s_LOGISIM_NET_313));

   NOT_GATE      GATE_130 (.Input_1(s_LOGISIM_NET_7),
                           .Result(s_LOGISIM_NET_273));

   AND_GATE_7_INPUTS #(.BubblesMask(0))
      GATE_131 (.Input_1(s_LOGISIM_NET_155),
                .Input_2(s_LOGISIM_NET_256),
                .Input_3(s_LOGISIM_NET_9),
                .Input_4(s_LOGISIM_NET_396),
                .Input_5(s_LOGISIM_NET_265),
                .Input_6(s_LOGISIM_NET_7),
                .Input_7(s_LOGISIM_NET_5),
                .Result(s_LOGISIM_NET_335));

   NOT_GATE      GATE_132 (.Input_1(s_LOGISIM_NET_22),
                           .Result(s_LOGISIM_NET_314));

   NOT_GATE      GATE_133 (.Input_1(s_LOGISIM_NET_22),
                           .Result(s_LOGISIM_NET_272));

   AND_GATE_10_INPUTS #(.BubblesMask(0))
      GATE_134 (.Input_1(s_LOGISIM_NET_286),
                .Input_10(s_LOGISIM_NET_18),
                .Input_2(s_LOGISIM_NET_227),
                .Input_3(s_LOGISIM_NET_9),
                .Input_4(s_LOGISIM_NET_32),
                .Input_5(s_LOGISIM_NET_147),
                .Input_6(s_LOGISIM_NET_35),
                .Input_7(s_LOGISIM_NET_48),
                .Input_8(s_LOGISIM_NET_5),
                .Input_9(s_LOGISIM_NET_53),
                .Result(s_LOGISIM_NET_257));

   NOT_GATE      GATE_135 (.Input_1(s_LOGISIM_NET_5),
                           .Result(s_LOGISIM_NET_276));

   NOT_GATE      GATE_136 (.Input_1(s_LOGISIM_NET_10),
                           .Result(s_LOGISIM_NET_277));

   NOT_GATE      GATE_137 (.Input_1(s_LOGISIM_NET_10),
                           .Result(s_LOGISIM_NET_221));

   NOT_GATE      GATE_138 (.Input_1(s_LOGISIM_NET_35),
                           .Result(s_LOGISIM_NET_400));

   NOT_GATE      GATE_139 (.Input_1(s_LOGISIM_NET_31),
                           .Result(s_LOGISIM_NET_40));

   NOT_GATE      GATE_140 (.Input_1(s_LOGISIM_NET_32),
                           .Result(s_LOGISIM_NET_27));

   NOT_GATE      GATE_141 (.Input_1(s_LOGISIM_NET_5),
                           .Result(s_LOGISIM_NET_310));

   NOT_GATE      GATE_142 (.Input_1(s_LOGISIM_NET_7),
                           .Result(s_LOGISIM_NET_48));

   NOT_GATE      GATE_143 (.Input_1(s_LOGISIM_NET_14),
                           .Result(s_LOGISIM_NET_143));

   NOT_GATE      GATE_144 (.Input_1(s_LOGISIM_NET_35),
                           .Result(s_LOGISIM_NET_102));

   NOT_GATE      GATE_145 (.Input_1(s_LOGISIM_NET_14),
                           .Result(s_LOGISIM_NET_332));

   NOT_GATE      GATE_146 (.Input_1(s_LOGISIM_NET_31),
                           .Result(s_LOGISIM_NET_88));

   NOT_GATE      GATE_147 (.Input_1(s_LOGISIM_NET_10),
                           .Result(s_LOGISIM_NET_154));

   NOT_GATE      GATE_148 (.Input_1(s_LOGISIM_NET_14),
                           .Result(s_LOGISIM_NET_20));

   NOT_GATE      GATE_149 (.Input_1(s_LOGISIM_NET_7),
                           .Result(s_LOGISIM_NET_172));

   NOT_GATE      GATE_150 (.Input_1(s_LOGISIM_NET_35),
                           .Result(s_LOGISIM_NET_94));

   NOT_GATE      GATE_151 (.Input_1(s_LOGISIM_NET_9),
                           .Result(s_LOGISIM_NET_362));

   NOT_GATE      GATE_152 (.Input_1(s_LOGISIM_NET_22),
                           .Result(s_LOGISIM_NET_137));

   NOT_GATE      GATE_153 (.Input_1(s_LOGISIM_NET_9),
                           .Result(s_LOGISIM_NET_186));

   NOT_GATE      GATE_154 (.Input_1(s_LOGISIM_NET_14),
                           .Result(s_LOGISIM_NET_111));

   NOT_GATE      GATE_155 (.Input_1(s_LOGISIM_NET_10),
                           .Result(s_LOGISIM_NET_352));

   NOT_GATE      GATE_156 (.Input_1(s_LOGISIM_NET_14),
                           .Result(s_LOGISIM_NET_303));

   NOT_GATE      GATE_157 (.Input_1(s_LOGISIM_NET_31),
                           .Result(s_LOGISIM_NET_47));

   NOT_GATE      GATE_158 (.Input_1(s_LOGISIM_NET_22),
                           .Result(s_LOGISIM_NET_179));

   NOT_GATE      GATE_159 (.Input_1(s_LOGISIM_NET_22),
                           .Result(s_LOGISIM_NET_39));

   AND_GATE_10_INPUTS #(.BubblesMask(0))
      GATE_160 (.Input_1(s_LOGISIM_NET_18),
                .Input_10(s_LOGISIM_NET_20),
                .Input_2(s_LOGISIM_NET_234),
                .Input_3(s_LOGISIM_NET_5),
                .Input_4(s_LOGISIM_NET_185),
                .Input_5(s_LOGISIM_NET_35),
                .Input_6(s_LOGISIM_NET_299),
                .Input_7(s_LOGISIM_NET_139),
                .Input_8(s_LOGISIM_NET_9),
                .Input_9(s_LOGISIM_NET_146),
                .Result(s_LOGISIM_NET_331));

   NOT_GATE      GATE_161 (.Input_1(s_LOGISIM_NET_31),
                           .Result(s_LOGISIM_NET_355));

   NOT_GATE      GATE_162 (.Input_1(s_LOGISIM_NET_35),
                           .Result(s_LOGISIM_NET_309));

   NOT_GATE      GATE_163 (.Input_1(s_LOGISIM_NET_14),
                           .Result(s_LOGISIM_NET_100));

   NOT_GATE      GATE_164 (.Input_1(s_LOGISIM_NET_7),
                           .Result(s_LOGISIM_NET_181));

   NOT_GATE      GATE_165 (.Input_1(s_LOGISIM_NET_32),
                           .Result(s_LOGISIM_NET_368));

   AND_GATE_7_INPUTS #(.BubblesMask(0))
      GATE_166 (.Input_1(s_LOGISIM_NET_135),
                .Input_2(s_LOGISIM_NET_247),
                .Input_3(s_LOGISIM_NET_32),
                .Input_4(s_LOGISIM_NET_31),
                .Input_5(s_LOGISIM_NET_202),
                .Input_6(s_LOGISIM_NET_379),
                .Input_7(s_LOGISIM_NET_205),
                .Result(s_LOGISIM_NET_217));

   NOT_GATE      GATE_167 (.Input_1(s_LOGISIM_NET_22),
                           .Result(s_LOGISIM_NET_157));

   NOT_GATE      GATE_168 (.Input_1(s_LOGISIM_NET_35),
                           .Result(s_LOGISIM_NET_178));

   NOT_GATE      GATE_169 (.Input_1(s_LOGISIM_NET_18),
                           .Result(s_LOGISIM_NET_237));

   AND_GATE_10_INPUTS #(.BubblesMask(0))
      GATE_170 (.Input_1(s_LOGISIM_NET_189),
                .Input_10(s_LOGISIM_NET_149),
                .Input_2(s_LOGISIM_NET_221),
                .Input_3(s_LOGISIM_NET_78),
                .Input_4(s_LOGISIM_NET_301),
                .Input_5(s_LOGISIM_NET_316),
                .Input_6(s_LOGISIM_NET_198),
                .Input_7(s_LOGISIM_NET_32),
                .Input_8(s_LOGISIM_NET_9),
                .Input_9(s_LOGISIM_NET_270),
                .Result(s_LOGISIM_NET_293));

   NOT_GATE      GATE_171 (.Input_1(s_LOGISIM_NET_32),
                           .Result(s_LOGISIM_NET_393));

   AND_GATE_7_INPUTS #(.BubblesMask(0))
      GATE_172 (.Input_1(s_LOGISIM_NET_42),
                .Input_2(s_LOGISIM_NET_197),
                .Input_3(s_LOGISIM_NET_9),
                .Input_4(s_LOGISIM_NET_267),
                .Input_5(s_LOGISIM_NET_103),
                .Input_6(s_LOGISIM_NET_5),
                .Input_7(s_LOGISIM_NET_380),
                .Result(s_LOGISIM_NET_3));

   NOT_GATE      GATE_173 (.Input_1(s_LOGISIM_NET_35),
                           .Result(s_LOGISIM_NET_321));

   AND_GATE_9_INPUTS #(.BubblesMask(0))
      GATE_174 (.Input_1(s_LOGISIM_NET_216),
                .Input_2(s_LOGISIM_NET_137),
                .Input_3(s_LOGISIM_NET_9),
                .Input_4(s_LOGISIM_NET_246),
                .Input_5(s_LOGISIM_NET_35),
                .Input_6(s_LOGISIM_NET_203),
                .Input_7(s_LOGISIM_NET_5),
                .Input_8(s_LOGISIM_NET_82),
                .Input_9(s_LOGISIM_NET_18),
                .Result(s_LOGISIM_NET_44));

   NOT_GATE      GATE_175 (.Input_1(s_LOGISIM_NET_14),
                           .Result(s_LOGISIM_NET_52));

   AND_GATE_6_INPUTS #(.BubblesMask(0))
      GATE_176 (.Input_1(s_LOGISIM_NET_72),
                .Input_2(s_LOGISIM_NET_170),
                .Input_3(s_LOGISIM_NET_9),
                .Input_4(s_LOGISIM_NET_283),
                .Input_5(s_LOGISIM_NET_226),
                .Input_6(s_LOGISIM_NET_375),
                .Result(s_LOGISIM_NET_104));

   NOT_GATE      GATE_177 (.Input_1(s_LOGISIM_NET_31),
                           .Result(s_LOGISIM_NET_350));

   AND_GATE_8_INPUTS #(.BubblesMask(0))
      GATE_178 (.Input_1(s_LOGISIM_NET_105),
                .Input_2(s_LOGISIM_NET_248),
                .Input_3(s_LOGISIM_NET_9),
                .Input_4(s_LOGISIM_NET_79),
                .Input_5(s_LOGISIM_NET_342),
                .Input_6(s_LOGISIM_NET_54),
                .Input_7(s_LOGISIM_NET_345),
                .Input_8(s_LOGISIM_NET_67),
                .Result(s_LOGISIM_NET_295));

   NOT_GATE      GATE_179 (.Input_1(s_LOGISIM_NET_22),
                           .Result(s_LOGISIM_NET_74));

   NOT_GATE      GATE_180 (.Input_1(s_LOGISIM_NET_7),
                           .Result(s_LOGISIM_NET_50));

   NOT_GATE      GATE_181 (.Input_1(s_LOGISIM_NET_10),
                           .Result(s_LOGISIM_NET_141));

   NOT_GATE      GATE_182 (.Input_1(s_LOGISIM_NET_22),
                           .Result(s_LOGISIM_NET_253));

   NOT_GATE      GATE_183 (.Input_1(s_LOGISIM_NET_7),
                           .Result(s_LOGISIM_NET_230));

   NOT_GATE      GATE_184 (.Input_1(s_LOGISIM_NET_31),
                           .Result(s_LOGISIM_NET_63));

   NOT_GATE      GATE_185 (.Input_1(s_LOGISIM_NET_35),
                           .Result(s_LOGISIM_NET_55));

   NOT_GATE      GATE_186 (.Input_1(s_LOGISIM_NET_14),
                           .Result(s_LOGISIM_NET_187));

   NOT_GATE      GATE_187 (.Input_1(s_LOGISIM_NET_9),
                           .Result(s_LOGISIM_NET_167));

   NOT_GATE      GATE_188 (.Input_1(s_LOGISIM_NET_14),
                           .Result(s_LOGISIM_NET_125));

   NOT_GATE      GATE_189 (.Input_1(s_LOGISIM_NET_18),
                           .Result(s_LOGISIM_NET_58));

   NOT_GATE      GATE_190 (.Input_1(s_LOGISIM_NET_35),
                           .Result(s_LOGISIM_NET_292));

   NOT_GATE      GATE_191 (.Input_1(s_LOGISIM_NET_22),
                           .Result(s_LOGISIM_NET_336));

   NOT_GATE      GATE_192 (.Input_1(s_LOGISIM_NET_31),
                           .Result(s_LOGISIM_NET_103));

   NOT_GATE      GATE_193 (.Input_1(s_LOGISIM_NET_5),
                           .Result(s_LOGISIM_NET_225));

   NOT_GATE      GATE_194 (.Input_1(s_LOGISIM_NET_7),
                           .Result(s_LOGISIM_NET_341));

   NOT_GATE      GATE_195 (.Input_1(s_LOGISIM_NET_14),
                           .Result(s_LOGISIM_NET_156));

   NOT_GATE      GATE_196 (.Input_1(s_LOGISIM_NET_18),
                           .Result(s_LOGISIM_NET_64));

   NOT_GATE      GATE_197 (.Input_1(s_LOGISIM_NET_31),
                           .Result(s_LOGISIM_NET_294));

   NOT_GATE      GATE_198 (.Input_1(s_LOGISIM_NET_18),
                           .Result(s_LOGISIM_NET_75));

   AND_GATE_10_INPUTS #(.BubblesMask(0))
      GATE_199 (.Input_1(s_LOGISIM_NET_18),
                .Input_10(s_LOGISIM_NET_111),
                .Input_2(s_LOGISIM_NET_1),
                .Input_3(s_LOGISIM_NET_5),
                .Input_4(s_LOGISIM_NET_168),
                .Input_5(s_LOGISIM_NET_35),
                .Input_6(s_LOGISIM_NET_397),
                .Input_7(s_LOGISIM_NET_32),
                .Input_8(s_LOGISIM_NET_9),
                .Input_9(s_LOGISIM_NET_24),
                .Result(s_LOGISIM_NET_131));

   NOT_GATE      GATE_200 (.Input_1(s_LOGISIM_NET_14),
                           .Result(s_LOGISIM_NET_15));

   NOT_GATE      GATE_201 (.Input_1(s_LOGISIM_NET_22),
                           .Result(s_LOGISIM_NET_33));

   NOT_GATE      GATE_202 (.Input_1(s_LOGISIM_NET_35),
                           .Result(s_LOGISIM_NET_316));

   NOT_GATE      GATE_203 (.Input_1(s_LOGISIM_NET_32),
                           .Result(s_LOGISIM_NET_267));

   NOT_GATE      GATE_204 (.Input_1(s_LOGISIM_NET_9),
                           .Result(s_LOGISIM_NET_30));

   NOT_GATE      GATE_205 (.Input_1(s_LOGISIM_NET_7),
                           .Result(s_LOGISIM_NET_43));

   NOT_GATE      GATE_206 (.Input_1(s_LOGISIM_NET_22),
                           .Result(s_LOGISIM_NET_146));

   NOT_GATE      GATE_207 (.Input_1(s_LOGISIM_NET_22),
                           .Result(s_LOGISIM_NET_196));

   NOT_GATE      GATE_208 (.Input_1(s_LOGISIM_NET_35),
                           .Result(s_LOGISIM_NET_11));

   NOT_GATE      GATE_209 (.Input_1(s_LOGISIM_NET_22),
                           .Result(s_LOGISIM_NET_197));

   NOT_GATE      GATE_210 (.Input_1(s_LOGISIM_NET_22),
                           .Result(s_LOGISIM_NET_306));

   NOT_GATE      GATE_211 (.Input_1(s_LOGISIM_NET_35),
                           .Result(s_LOGISIM_NET_202));

   AND_GATE_5_INPUTS #(.BubblesMask(0))
      GATE_212 (.Input_1(s_LOGISIM_NET_31),
                .Input_2(s_LOGISIM_NET_32),
                .Input_3(s_LOGISIM_NET_261),
                .Input_4(s_LOGISIM_NET_22),
                .Input_5(s_LOGISIM_NET_14),
                .Result(s_LOGISIM_NET_66));

   NOT_GATE      GATE_213 (.Input_1(s_LOGISIM_NET_32),
                           .Result(s_LOGISIM_NET_151));

   NOT_GATE      GATE_214 (.Input_1(s_LOGISIM_NET_35),
                           .Result(s_LOGISIM_NET_317));

   NOT_GATE      GATE_215 (.Input_1(s_LOGISIM_NET_5),
                           .Result(s_LOGISIM_NET_363));

   NOT_GATE      GATE_216 (.Input_1(s_LOGISIM_NET_32),
                           .Result(s_LOGISIM_NET_324));

   NOT_GATE      GATE_217 (.Input_1(s_LOGISIM_NET_35),
                           .Result(s_LOGISIM_NET_326));

   NOT_GATE      GATE_218 (.Input_1(s_LOGISIM_NET_22),
                           .Result(s_LOGISIM_NET_275));

   NOT_GATE      GATE_219 (.Input_1(s_LOGISIM_NET_5),
                           .Result(s_LOGISIM_NET_162));

   NOT_GATE      GATE_220 (.Input_1(s_LOGISIM_NET_35),
                           .Result(s_LOGISIM_NET_83));

   AND_GATE_7_INPUTS #(.BubblesMask(0))
      GATE_221 (.Input_1(s_LOGISIM_NET_281),
                .Input_2(s_LOGISIM_NET_126),
                .Input_3(s_LOGISIM_NET_9),
                .Input_4(s_LOGISIM_NET_368),
                .Input_5(s_LOGISIM_NET_136),
                .Input_6(s_LOGISIM_NET_7),
                .Input_7(s_LOGISIM_NET_5),
                .Result(s_LOGISIM_NET_207));

   NOT_GATE      GATE_222 (.Input_1(s_LOGISIM_NET_31),
                           .Result(s_LOGISIM_NET_349));

   NOT_GATE      GATE_223 (.Input_1(s_LOGISIM_NET_14),
                           .Result(s_LOGISIM_NET_255));

   NOT_GATE      GATE_224 (.Input_1(s_LOGISIM_NET_10),
                           .Result(s_LOGISIM_NET_12));

   NOT_GATE      GATE_225 (.Input_1(s_LOGISIM_NET_35),
                           .Result(s_LOGISIM_NET_245));

   NOT_GATE      GATE_226 (.Input_1(s_LOGISIM_NET_22),
                           .Result(s_LOGISIM_NET_365));

   NOT_GATE      GATE_227 (.Input_1(s_LOGISIM_NET_7),
                           .Result(s_LOGISIM_NET_108));

   AND_GATE_8_INPUTS #(.BubblesMask(0))
      GATE_228 (.Input_1(s_LOGISIM_NET_25),
                .Input_2(s_LOGISIM_NET_39),
                .Input_3(s_LOGISIM_NET_274),
                .Input_4(s_LOGISIM_NET_32),
                .Input_5(s_LOGISIM_NET_31),
                .Input_6(s_LOGISIM_NET_35),
                .Input_7(s_LOGISIM_NET_231),
                .Input_8(s_LOGISIM_NET_232),
                .Result(s_LOGISIM_NET_2));

   AND_GATE_8_INPUTS #(.BubblesMask(0))
      GATE_229 (.Input_1(s_LOGISIM_NET_255),
                .Input_2(s_LOGISIM_NET_60),
                .Input_3(s_LOGISIM_NET_236),
                .Input_4(s_LOGISIM_NET_393),
                .Input_5(s_LOGISIM_NET_241),
                .Input_6(s_LOGISIM_NET_94),
                .Input_7(s_LOGISIM_NET_242),
                .Input_8(s_LOGISIM_NET_5),
                .Result(s_LOGISIM_NET_26));

   NOT_GATE      GATE_230 (.Input_1(s_LOGISIM_NET_7),
                           .Result(s_LOGISIM_NET_168));

   NOT_GATE      GATE_231 (.Input_1(s_LOGISIM_NET_35),
                           .Result(s_LOGISIM_NET_360));

   NOT_GATE      GATE_232 (.Input_1(s_LOGISIM_NET_31),
                           .Result(s_LOGISIM_NET_300));

   AND_GATE_5_INPUTS #(.BubblesMask(0))
      GATE_233 (.Input_1(s_LOGISIM_NET_14),
                .Input_2(s_LOGISIM_NET_22),
                .Input_3(s_LOGISIM_NET_153),
                .Input_4(s_LOGISIM_NET_32),
                .Input_5(s_LOGISIM_NET_31),
                .Result(s_LOGISIM_NET_381));

   AND_GATE_8_INPUTS #(.BubblesMask(0))
      GATE_234 (.Input_1(s_LOGISIM_NET_276),
                .Input_2(s_LOGISIM_NET_7),
                .Input_3(s_LOGISIM_NET_228),
                .Input_4(s_LOGISIM_NET_250),
                .Input_5(s_LOGISIM_NET_151),
                .Input_6(s_LOGISIM_NET_235),
                .Input_7(s_LOGISIM_NET_387),
                .Input_8(s_LOGISIM_NET_92),
                .Result(s_LOGISIM_NET_318));

   NOT_GATE      GATE_235 (.Input_1(s_LOGISIM_NET_35),
                           .Result(s_LOGISIM_NET_132));

   NOT_GATE      GATE_236 (.Input_1(s_LOGISIM_NET_14),
                           .Result(s_LOGISIM_NET_149));

   NOT_GATE      GATE_237 (.Input_1(s_LOGISIM_NET_5),
                           .Result(s_LOGISIM_NET_232));

   NOT_GATE      GATE_238 (.Input_1(s_LOGISIM_NET_31),
                           .Result(s_LOGISIM_NET_390));

   NOT_GATE      GATE_239 (.Input_1(s_LOGISIM_NET_31),
                           .Result(s_LOGISIM_NET_391));

   NOT_GATE      GATE_240 (.Input_1(s_LOGISIM_NET_14),
                           .Result(s_LOGISIM_NET_174));

   AND_GATE_10_INPUTS #(.BubblesMask(0))
      GATE_241 (.Input_1(s_LOGISIM_NET_38),
                .Input_10(s_LOGISIM_NET_370),
                .Input_2(s_LOGISIM_NET_252),
                .Input_3(s_LOGISIM_NET_120),
                .Input_4(s_LOGISIM_NET_7),
                .Input_5(s_LOGISIM_NET_35),
                .Input_6(s_LOGISIM_NET_307),
                .Input_7(s_LOGISIM_NET_32),
                .Input_8(s_LOGISIM_NET_9),
                .Input_9(s_LOGISIM_NET_166),
                .Result(s_LOGISIM_NET_133));

   NOT_GATE      GATE_242 (.Input_1(s_LOGISIM_NET_35),
                           .Result(s_LOGISIM_NET_375));

   NOT_GATE      GATE_243 (.Input_1(s_LOGISIM_NET_22),
                           .Result(s_LOGISIM_NET_270));

   NOT_GATE      GATE_244 (.Input_1(s_LOGISIM_NET_5),
                           .Result(s_LOGISIM_NET_148));

   NOT_GATE      GATE_245 (.Input_1(s_LOGISIM_NET_7),
                           .Result(s_LOGISIM_NET_240));

   NOT_GATE      GATE_246 (.Input_1(s_LOGISIM_NET_7),
                           .Result(s_LOGISIM_NET_220));

   NOT_GATE      GATE_247 (.Input_1(s_LOGISIM_NET_7),
                           .Result(s_LOGISIM_NET_353));

   NOT_GATE      GATE_248 (.Input_1(s_LOGISIM_NET_31),
                           .Result(s_LOGISIM_NET_198));

   NOT_GATE      GATE_249 (.Input_1(s_LOGISIM_NET_5),
                           .Result(s_LOGISIM_NET_70));

   AND_GATE_7_INPUTS #(.BubblesMask(0))
      GATE_250 (.Input_1(s_LOGISIM_NET_322),
                .Input_2(s_LOGISIM_NET_183),
                .Input_3(s_LOGISIM_NET_343),
                .Input_4(s_LOGISIM_NET_32),
                .Input_5(s_LOGISIM_NET_31),
                .Input_6(s_LOGISIM_NET_230),
                .Input_7(s_LOGISIM_NET_363),
                .Result(s_LOGISIM_NET_269));

   NOT_GATE      GATE_251 (.Input_1(s_LOGISIM_NET_31),
                           .Result(s_LOGISIM_NET_291));

   NOT_GATE      GATE_252 (.Input_1(s_LOGISIM_NET_7),
                           .Result(s_LOGISIM_NET_330));

   AND_GATE_8_INPUTS #(.BubblesMask(0))
      GATE_253 (.Input_1(s_LOGISIM_NET_358),
                .Input_2(s_LOGISIM_NET_4),
                .Input_3(s_LOGISIM_NET_9),
                .Input_4(s_LOGISIM_NET_32),
                .Input_5(s_LOGISIM_NET_31),
                .Input_6(s_LOGISIM_NET_317),
                .Input_7(s_LOGISIM_NET_7),
                .Input_8(s_LOGISIM_NET_5),
                .Result(s_LOGISIM_NET_373));

   NOT_GATE      GATE_254 (.Input_1(s_LOGISIM_NET_9),
                           .Result(s_LOGISIM_NET_261));

   NOT_GATE      GATE_255 (.Input_1(s_LOGISIM_NET_9),
                           .Result(s_LOGISIM_NET_124));

   NOT_GATE      GATE_256 (.Input_1(s_LOGISIM_NET_5),
                           .Result(s_LOGISIM_NET_56));

   NOT_GATE      GATE_257 (.Input_1(s_LOGISIM_NET_22),
                           .Result(s_LOGISIM_NET_297));

   OR_GATE #(.BubblesMask(0))
      GATE_258 (.Input_1(s_LOGISIM_NET_128),
                .Input_2(s_LOGISIM_NET_388),
                .Result(s_LOGISIM_NET_377));

   NOT_GATE      GATE_259 (.Input_1(s_LOGISIM_NET_22),
                           .Result(s_LOGISIM_NET_117));

   AND_GATE_8_INPUTS #(.BubblesMask(0))
      GATE_260 (.Input_1(s_LOGISIM_NET_23),
                .Input_2(s_LOGISIM_NET_176),
                .Input_3(s_LOGISIM_NET_9),
                .Input_4(s_LOGISIM_NET_32),
                .Input_5(s_LOGISIM_NET_31),
                .Input_6(s_LOGISIM_NET_35),
                .Input_7(s_LOGISIM_NET_7),
                .Input_8(s_LOGISIM_NET_5),
                .Result(s_LOGISIM_NET_394));

   NOT_GATE      GATE_261 (.Input_1(s_LOGISIM_NET_7),
                           .Result(s_LOGISIM_NET_379));

   NOT_GATE      GATE_262 (.Input_1(s_LOGISIM_NET_5),
                           .Result(s_LOGISIM_NET_200));

   AND_GATE_7_INPUTS #(.BubblesMask(0))
      GATE_263 (.Input_1(s_LOGISIM_NET_125),
                .Input_2(s_LOGISIM_NET_280),
                .Input_3(s_LOGISIM_NET_194),
                .Input_4(s_LOGISIM_NET_32),
                .Input_5(s_LOGISIM_NET_31),
                .Input_6(s_LOGISIM_NET_171),
                .Input_7(s_LOGISIM_NET_243),
                .Result(s_LOGISIM_NET_348));

   NOT_GATE      GATE_264 (.Input_1(s_LOGISIM_NET_22),
                           .Result(s_LOGISIM_NET_6));

   NOT_GATE      GATE_265 (.Input_1(s_LOGISIM_NET_22),
                           .Result(s_LOGISIM_NET_287));

   NOT_GATE      GATE_266 (.Input_1(s_LOGISIM_NET_14),
                           .Result(s_LOGISIM_NET_358));

   NOT_GATE      GATE_267 (.Input_1(s_LOGISIM_NET_14),
                           .Result(s_LOGISIM_NET_155));

   NOT_GATE      GATE_268 (.Input_1(s_LOGISIM_NET_7),
                           .Result(s_LOGISIM_NET_374));

   NOT_GATE      GATE_269 (.Input_1(s_LOGISIM_NET_14),
                           .Result(s_LOGISIM_NET_99));

   NOT_GATE      GATE_270 (.Input_1(s_LOGISIM_NET_31),
                           .Result(s_LOGISIM_NET_327));

   NOT_GATE      GATE_271 (.Input_1(s_LOGISIM_NET_9),
                           .Result(s_LOGISIM_NET_153));

   NOT_GATE      GATE_272 (.Input_1(s_LOGISIM_NET_7),
                           .Result(s_LOGISIM_NET_242));

   NOT_GATE      GATE_273 (.Input_1(s_LOGISIM_NET_22),
                           .Result(s_LOGISIM_NET_227));

   NOT_GATE      GATE_274 (.Input_1(s_LOGISIM_NET_9),
                           .Result(s_LOGISIM_NET_49));

   NOT_GATE      GATE_275 (.Input_1(s_LOGISIM_NET_9),
                           .Result(s_LOGISIM_NET_93));

   AND_GATE_6_INPUTS #(.BubblesMask(0))
      GATE_276 (.Input_1(s_LOGISIM_NET_208),
                .Input_2(s_LOGISIM_NET_365),
                .Input_3(s_LOGISIM_NET_9),
                .Input_4(s_LOGISIM_NET_163),
                .Input_5(s_LOGISIM_NET_73),
                .Input_6(s_LOGISIM_NET_329),
                .Result(s_LOGISIM_NET_46));

   AND_GATE_10_INPUTS #(.BubblesMask(0))
      GATE_277 (.Input_1(s_LOGISIM_NET_222),
                .Input_10(s_LOGISIM_NET_282),
                .Input_2(s_LOGISIM_NET_154),
                .Input_3(s_LOGISIM_NET_5),
                .Input_4(s_LOGISIM_NET_7),
                .Input_5(s_LOGISIM_NET_35),
                .Input_6(s_LOGISIM_NET_113),
                .Input_7(s_LOGISIM_NET_32),
                .Input_8(s_LOGISIM_NET_9),
                .Input_9(s_LOGISIM_NET_84),
                .Result(s_LOGISIM_NET_211));

   NOT_GATE      GATE_278 (.Input_1(s_LOGISIM_NET_35),
                           .Result(s_LOGISIM_NET_182));

   NOT_GATE      GATE_279 (.Input_1(s_LOGISIM_NET_32),
                           .Result(s_LOGISIM_NET_173));

   NOT_GATE      GATE_280 (.Input_1(s_LOGISIM_NET_14),
                           .Result(s_LOGISIM_NET_90));

   NOT_GATE      GATE_281 (.Input_1(s_LOGISIM_NET_7),
                           .Result(s_LOGISIM_NET_320));

   NOT_GATE      GATE_282 (.Input_1(s_LOGISIM_NET_5),
                           .Result(s_LOGISIM_NET_213));

   NOT_GATE      GATE_283 (.Input_1(s_LOGISIM_NET_10),
                           .Result(s_LOGISIM_NET_252));

   NOT_GATE      GATE_284 (.Input_1(s_LOGISIM_NET_14),
                           .Result(s_LOGISIM_NET_77));

   NOT_GATE      GATE_285 (.Input_1(s_LOGISIM_NET_32),
                           .Result(s_LOGISIM_NET_346));

   NOT_GATE      GATE_286 (.Input_1(s_LOGISIM_NET_14),
                           .Result(s_LOGISIM_NET_96));

   NOT_GATE      GATE_287 (.Input_1(s_LOGISIM_NET_32),
                           .Result(s_LOGISIM_NET_79));

   NOT_GATE      GATE_288 (.Input_1(s_LOGISIM_NET_14),
                           .Result(s_LOGISIM_NET_72));

   NOT_GATE      GATE_289 (.Input_1(s_LOGISIM_NET_31),
                           .Result(s_LOGISIM_NET_210));

   NOT_GATE      GATE_290 (.Input_1(s_LOGISIM_NET_31),
                           .Result(s_LOGISIM_NET_342));

   NOT_GATE      GATE_291 (.Input_1(s_LOGISIM_NET_22),
                           .Result(s_LOGISIM_NET_161));

   NOT_GATE      GATE_292 (.Input_1(s_LOGISIM_NET_18),
                           .Result(s_LOGISIM_NET_304));

   NOT_GATE      GATE_293 (.Input_1(s_LOGISIM_NET_31),
                           .Result(s_LOGISIM_NET_285));

   AND_GATE_8_INPUTS #(.BubblesMask(0))
      GATE_294 (.Input_1(s_LOGISIM_NET_96),
                .Input_2(s_LOGISIM_NET_287),
                .Input_3(s_LOGISIM_NET_142),
                .Input_4(s_LOGISIM_NET_32),
                .Input_5(s_LOGISIM_NET_384),
                .Input_6(s_LOGISIM_NET_354),
                .Input_7(s_LOGISIM_NET_7),
                .Input_8(s_LOGISIM_NET_152),
                .Result(s_LOGISIM_NET_392));

   NOT_GATE      GATE_295 (.Input_1(s_LOGISIM_NET_14),
                           .Result(s_LOGISIM_NET_259));

   NOT_GATE      GATE_296 (.Input_1(s_LOGISIM_NET_14),
                           .Result(s_LOGISIM_NET_19));

   AND_GATE_8_INPUTS #(.BubblesMask(0))
      GATE_297 (.Input_1(s_LOGISIM_NET_5),
                .Input_2(s_LOGISIM_NET_220),
                .Input_3(s_LOGISIM_NET_11),
                .Input_4(s_LOGISIM_NET_349),
                .Input_5(s_LOGISIM_NET_27),
                .Input_6(s_LOGISIM_NET_9),
                .Input_7(s_LOGISIM_NET_33),
                .Input_8(s_LOGISIM_NET_174),
                .Result(s_LOGISIM_NET_191));

   NOT_GATE      GATE_298 (.Input_1(s_LOGISIM_NET_31),
                           .Result(s_LOGISIM_NET_241));

   NOT_GATE      GATE_299 (.Input_1(s_LOGISIM_NET_14),
                           .Result(s_LOGISIM_NET_298));

   NOT_GATE      GATE_300 (.Input_1(s_LOGISIM_NET_22),
                           .Result(s_LOGISIM_NET_206));

   NOT_GATE      GATE_301 (.Input_1(s_LOGISIM_NET_22),
                           .Result(s_LOGISIM_NET_170));

   NOT_GATE      GATE_302 (.Input_1(s_LOGISIM_NET_31),
                           .Result(s_LOGISIM_NET_218));

   NOT_GATE      GATE_303 (.Input_1(s_LOGISIM_NET_14),
                           .Result(s_LOGISIM_NET_322));

   NOT_GATE      GATE_304 (.Input_1(s_LOGISIM_NET_22),
                           .Result(s_LOGISIM_NET_123));

   OR_GATE_6_INPUTS #(.BubblesMask(0))
      GATE_305 (.Input_1(s_LOGISIM_NET_138),
                .Input_2(s_LOGISIM_NET_348),
                .Input_3(s_LOGISIM_NET_269),
                .Input_4(s_LOGISIM_NET_127),
                .Input_5(s_LOGISIM_NET_385),
                .Input_6(s_LOGISIM_NET_257),
                .Result(s_LOGISIM_NET_383));

   NOT_GATE      GATE_306 (.Input_1(s_LOGISIM_NET_22),
                           .Result(s_LOGISIM_NET_256));

   NOT_GATE      GATE_307 (.Input_1(s_LOGISIM_NET_18),
                           .Result(s_LOGISIM_NET_150));

   NOT_GATE      GATE_308 (.Input_1(s_LOGISIM_NET_9),
                           .Result(s_LOGISIM_NET_107));

   NOT_GATE      GATE_309 (.Input_1(s_LOGISIM_NET_10),
                           .Result(s_LOGISIM_NET_82));

   NOT_GATE      GATE_310 (.Input_1(s_LOGISIM_NET_5),
                           .Result(s_LOGISIM_NET_271));

   OR_GATE_21_INPUTS #(.BubblesMask(0))
      GATE_311 (.Input_1(s_LOGISIM_NET_293),
                .Input_10(s_LOGISIM_NET_191),
                .Input_11(s_LOGISIM_NET_398),
                .Input_12(s_LOGISIM_NET_366),
                .Input_13(s_LOGISIM_NET_69),
                .Input_14(s_LOGISIM_NET_331),
                .Input_15(s_LOGISIM_NET_318),
                .Input_16(s_LOGISIM_NET_66),
                .Input_17(s_LOGISIM_NET_356),
                .Input_18(s_LOGISIM_NET_131),
                .Input_19(s_LOGISIM_NET_361),
                .Input_2(s_LOGISIM_NET_85),
                .Input_20(s_LOGISIM_NET_41),
                .Input_21(s_LOGISIM_NET_34),
                .Input_3(s_LOGISIM_NET_211),
                .Input_4(s_LOGISIM_NET_91),
                .Input_5(s_LOGISIM_NET_116),
                .Input_6(s_LOGISIM_NET_133),
                .Input_7(s_LOGISIM_NET_239),
                .Input_8(s_LOGISIM_NET_17),
                .Input_9(s_LOGISIM_NET_112),
                .Result(s_LOGISIM_NET_389));

   NOT_GATE      GATE_312 (.Input_1(s_LOGISIM_NET_32),
                           .Result(s_LOGISIM_NET_262));

   AND_GATE_8_INPUTS #(.BubblesMask(0))
      GATE_313 (.Input_1(s_LOGISIM_NET_308),
                .Input_2(s_LOGISIM_NET_206),
                .Input_3(s_LOGISIM_NET_49),
                .Input_4(s_LOGISIM_NET_32),
                .Input_5(s_LOGISIM_NET_31),
                .Input_6(s_LOGISIM_NET_309),
                .Input_7(s_LOGISIM_NET_160),
                .Input_8(s_LOGISIM_NET_5),
                .Result(s_LOGISIM_NET_369));

   NOT_GATE      GATE_314 (.Input_1(s_LOGISIM_NET_9),
                           .Result(s_LOGISIM_NET_235));

   NOT_GATE      GATE_315 (.Input_1(s_LOGISIM_NET_5),
                           .Result(s_LOGISIM_NET_57));

   NOT_GATE      GATE_316 (.Input_1(s_LOGISIM_NET_35),
                           .Result(s_LOGISIM_NET_134));

   NOT_GATE      GATE_317 (.Input_1(s_LOGISIM_NET_14),
                           .Result(s_LOGISIM_NET_42));

   NOT_GATE      GATE_318 (.Input_1(s_LOGISIM_NET_22),
                           .Result(s_LOGISIM_NET_311));

   NOT_GATE      GATE_319 (.Input_1(s_LOGISIM_NET_10),
                           .Result(s_LOGISIM_NET_129));

   NOT_GATE      GATE_320 (.Input_1(s_LOGISIM_NET_5),
                           .Result(s_LOGISIM_NET_152));

   NOT_GATE      GATE_321 (.Input_1(s_LOGISIM_NET_7),
                           .Result(s_LOGISIM_NET_301));

   NOT_GATE      GATE_322 (.Input_1(s_LOGISIM_NET_22),
                           .Result(s_LOGISIM_NET_190));

   NOT_GATE      GATE_323 (.Input_1(s_LOGISIM_NET_31),
                           .Result(s_LOGISIM_NET_119));

   NOT_GATE      GATE_324 (.Input_1(s_LOGISIM_NET_14),
                           .Result(s_LOGISIM_NET_281));

   AND_GATE_10_INPUTS #(.BubblesMask(0))
      GATE_325 (.Input_1(s_LOGISIM_NET_209),
                .Input_10(s_LOGISIM_NET_15),
                .Input_2(s_LOGISIM_NET_315),
                .Input_3(s_LOGISIM_NET_213),
                .Input_4(s_LOGISIM_NET_7),
                .Input_5(s_LOGISIM_NET_326),
                .Input_6(s_LOGISIM_NET_218),
                .Input_7(s_LOGISIM_NET_32),
                .Input_8(s_LOGISIM_NET_9),
                .Input_9(s_LOGISIM_NET_288),
                .Result(s_LOGISIM_NET_116));

   NOT_GATE      GATE_326 (.Input_1(s_LOGISIM_NET_18),
                           .Result(s_LOGISIM_NET_38));

   NOT_GATE      GATE_327 (.Input_1(s_LOGISIM_NET_7),
                           .Result(s_LOGISIM_NET_36));

   NOT_GATE      GATE_328 (.Input_1(s_LOGISIM_NET_5),
                           .Result(s_LOGISIM_NET_205));

   NOT_GATE      GATE_329 (.Input_1(s_LOGISIM_NET_14),
                           .Result(s_LOGISIM_NET_101));

   AND_GATE_8_INPUTS #(.BubblesMask(0))
      GATE_330 (.Input_1(s_LOGISIM_NET_258),
                .Input_2(s_LOGISIM_NET_122),
                .Input_3(s_LOGISIM_NET_9),
                .Input_4(s_LOGISIM_NET_229),
                .Input_5(s_LOGISIM_NET_119),
                .Input_6(s_LOGISIM_NET_214),
                .Input_7(s_LOGISIM_NET_382),
                .Input_8(s_LOGISIM_NET_64),
                .Result(s_LOGISIM_NET_333));

   OR_GATE_11_INPUTS #(.BubblesMask(0))
      GATE_331 (.Input_1(s_LOGISIM_NET_164),
                .Input_10(s_LOGISIM_NET_44),
                .Input_11(s_LOGISIM_NET_251),
                .Input_2(s_LOGISIM_NET_323),
                .Input_3(s_LOGISIM_NET_177),
                .Input_4(s_LOGISIM_NET_158),
                .Input_5(s_LOGISIM_NET_217),
                .Input_6(s_LOGISIM_NET_46),
                .Input_7(s_LOGISIM_NET_295),
                .Input_8(s_LOGISIM_NET_204),
                .Input_9(s_LOGISIM_NET_335),
                .Result(s_LOGISIM_NET_372));

   NOT_GATE      GATE_332 (.Input_1(s_LOGISIM_NET_5),
                           .Result(s_LOGISIM_NET_114));

   NOT_GATE      GATE_333 (.Input_1(s_LOGISIM_NET_10),
                           .Result(s_LOGISIM_NET_263));

   NOT_GATE      GATE_334 (.Input_1(s_LOGISIM_NET_5),
                           .Result(s_LOGISIM_NET_254));

   NOT_GATE      GATE_335 (.Input_1(s_LOGISIM_NET_22),
                           .Result(s_LOGISIM_NET_126));

   NOT_GATE      GATE_336 (.Input_1(s_LOGISIM_NET_5),
                           .Result(s_LOGISIM_NET_347));

   AND_GATE_8_INPUTS #(.BubblesMask(0))
      GATE_337 (.Input_1(s_LOGISIM_NET_100),
                .Input_2(s_LOGISIM_NET_313),
                .Input_3(s_LOGISIM_NET_167),
                .Input_4(s_LOGISIM_NET_193),
                .Input_5(s_LOGISIM_NET_63),
                .Input_6(s_LOGISIM_NET_178),
                .Input_7(s_LOGISIM_NET_374),
                .Input_8(s_LOGISIM_NET_5),
                .Result(s_LOGISIM_NET_128));

   NOT_GATE      GATE_338 (.Input_1(s_LOGISIM_NET_14),
                           .Result(s_LOGISIM_NET_81));

   NOT_GATE      GATE_339 (.Input_1(s_LOGISIM_NET_31),
                           .Result(s_LOGISIM_NET_266));

   NOT_GATE      GATE_340 (.Input_1(s_LOGISIM_NET_10),
                           .Result(s_LOGISIM_NET_315));

   NOT_GATE      GATE_341 (.Input_1(s_LOGISIM_NET_9),
                           .Result(s_LOGISIM_NET_236));

   AND_GATE_7_INPUTS #(.BubblesMask(0))
      GATE_342 (.Input_1(s_LOGISIM_NET_180),
                .Input_2(s_LOGISIM_NET_275),
                .Input_3(s_LOGISIM_NET_186),
                .Input_4(s_LOGISIM_NET_47),
                .Input_5(s_LOGISIM_NET_338),
                .Input_6(s_LOGISIM_NET_7),
                .Input_7(s_LOGISIM_NET_310),
                .Result(s_LOGISIM_NET_290));

   NOT_GATE      GATE_343 (.Input_1(s_LOGISIM_NET_32),
                           .Result(s_LOGISIM_NET_139));

   AND_GATE_8_INPUTS #(.BubblesMask(0))
      GATE_344 (.Input_1(s_LOGISIM_NET_45),
                .Input_2(s_LOGISIM_NET_249),
                .Input_3(s_LOGISIM_NET_30),
                .Input_4(s_LOGISIM_NET_32),
                .Input_5(s_LOGISIM_NET_199),
                .Input_6(s_LOGISIM_NET_55),
                .Input_7(s_LOGISIM_NET_7),
                .Input_8(s_LOGISIM_NET_57),
                .Result(s_LOGISIM_NET_138));

   NOT_GATE      GATE_345 (.Input_1(s_LOGISIM_NET_14),
                           .Result(s_LOGISIM_NET_286));

   AND_GATE_8_INPUTS #(.BubblesMask(0))
      GATE_346 (.Input_1(s_LOGISIM_NET_81),
                .Input_2(s_LOGISIM_NET_157),
                .Input_3(s_LOGISIM_NET_296),
                .Input_4(s_LOGISIM_NET_402),
                .Input_5(s_LOGISIM_NET_302),
                .Input_6(s_LOGISIM_NET_97),
                .Input_7(s_LOGISIM_NET_7),
                .Input_8(s_LOGISIM_NET_59),
                .Result(s_LOGISIM_NET_388));

   NOT_GATE      GATE_347 (.Input_1(s_LOGISIM_NET_35),
                           .Result(s_LOGISIM_NET_260));

   NOT_GATE      GATE_348 (.Input_1(s_LOGISIM_NET_22),
                           .Result(s_LOGISIM_NET_279));

   NOT_GATE      GATE_349 (.Input_1(s_LOGISIM_NET_35),
                           .Result(s_LOGISIM_NET_329));

   NOT_GATE      GATE_350 (.Input_1(s_LOGISIM_NET_10),
                           .Result(s_LOGISIM_NET_234));

   NOT_GATE      GATE_351 (.Input_1(s_LOGISIM_NET_14),
                           .Result(s_LOGISIM_NET_105));

   NOT_GATE      GATE_352 (.Input_1(s_LOGISIM_NET_9),
                           .Result(s_LOGISIM_NET_247));

   NOT_GATE      GATE_353 (.Input_1(s_LOGISIM_NET_10),
                           .Result(s_LOGISIM_NET_53));

   AND_GATE_10_INPUTS #(.BubblesMask(0))
      GATE_354 (.Input_1(s_LOGISIM_NET_304),
                .Input_10(s_LOGISIM_NET_61),
                .Input_2(s_LOGISIM_NET_141),
                .Input_3(s_LOGISIM_NET_271),
                .Input_4(s_LOGISIM_NET_106),
                .Input_5(s_LOGISIM_NET_35),
                .Input_6(s_LOGISIM_NET_391),
                .Input_7(s_LOGISIM_NET_346),
                .Input_8(s_LOGISIM_NET_9),
                .Input_9(s_LOGISIM_NET_117),
                .Result(s_LOGISIM_NET_366));

   NOT_GATE      GATE_355 (.Input_1(s_LOGISIM_NET_35),
                           .Result(s_LOGISIM_NET_312));

   NOT_GATE      GATE_356 (.Input_1(s_LOGISIM_NET_32),
                           .Result(s_LOGISIM_NET_13));

   NOT_GATE      GATE_357 (.Input_1(s_LOGISIM_NET_14),
                           .Result(s_LOGISIM_NET_215));

   NOT_GATE      GATE_358 (.Input_1(s_LOGISIM_NET_14),
                           .Result(s_LOGISIM_NET_192));

   NOT_GATE      GATE_359 (.Input_1(s_LOGISIM_NET_10),
                           .Result(s_LOGISIM_NET_165));

   NOT_GATE      GATE_360 (.Input_1(s_LOGISIM_NET_14),
                           .Result(s_LOGISIM_NET_208));

   AND_GATE_5_INPUTS #(.BubblesMask(0))
      GATE_361 (.Input_1(s_LOGISIM_NET_14),
                .Input_2(s_LOGISIM_NET_367),
                .Input_3(s_LOGISIM_NET_9),
                .Input_4(s_LOGISIM_NET_109),
                .Input_5(s_LOGISIM_NET_294),
                .Result(s_LOGISIM_NET_401));

   NOT_GATE      GATE_362 (.Input_1(s_LOGISIM_NET_14),
                           .Result(s_LOGISIM_NET_180));

   NOT_GATE      GATE_363 (.Input_1(s_LOGISIM_NET_32),
                           .Result(s_LOGISIM_NET_283));

   NOT_GATE      GATE_364 (.Input_1(s_LOGISIM_NET_35),
                           .Result(s_LOGISIM_NET_201));

   NOT_GATE      GATE_365 (.Input_1(s_LOGISIM_NET_35),
                           .Result(s_LOGISIM_NET_97));

   NOT_GATE      GATE_366 (.Input_1(s_LOGISIM_NET_35),
                           .Result(s_LOGISIM_NET_354));

   NOT_GATE      GATE_367 (.Input_1(s_LOGISIM_NET_32),
                           .Result(s_LOGISIM_NET_65));

   NOT_GATE      GATE_368 (.Input_1(s_LOGISIM_NET_31),
                           .Result(s_LOGISIM_NET_136));

   AND_GATE_8_INPUTS #(.BubblesMask(0))
      GATE_369 (.Input_1(s_LOGISIM_NET_52),
                .Input_2(s_LOGISIM_NET_159),
                .Input_3(s_LOGISIM_NET_9),
                .Input_4(s_LOGISIM_NET_32),
                .Input_5(s_LOGISIM_NET_88),
                .Input_6(s_LOGISIM_NET_7),
                .Input_7(s_LOGISIM_NET_165),
                .Input_8(s_LOGISIM_NET_58),
                .Result(s_LOGISIM_NET_385));

   NOT_GATE      GATE_370 (.Input_1(s_LOGISIM_NET_31),
                           .Result(s_LOGISIM_NET_265));

   NOT_GATE      GATE_371 (.Input_1(s_LOGISIM_NET_22),
                           .Result(s_LOGISIM_NET_166));

   NOT_GATE      GATE_372 (.Input_1(s_LOGISIM_NET_22),
                           .Result(s_LOGISIM_NET_183));

   NOT_GATE      GATE_373 (.Input_1(s_LOGISIM_NET_22),
                           .Result(s_LOGISIM_NET_175));

   NOT_GATE      GATE_374 (.Input_1(s_LOGISIM_NET_18),
                           .Result(s_LOGISIM_NET_140));

   NOT_GATE      GATE_375 (.Input_1(s_LOGISIM_NET_22),
                           .Result(s_LOGISIM_NET_387));

   NOT_GATE      GATE_376 (.Input_1(s_LOGISIM_NET_22),
                           .Result(s_LOGISIM_NET_249));

   NOT_GATE      GATE_377 (.Input_1(s_LOGISIM_NET_10),
                           .Result(s_LOGISIM_NET_95));

   AND_GATE_8_INPUTS #(.BubblesMask(0))
      GATE_378 (.Input_1(s_LOGISIM_NET_200),
                .Input_2(s_LOGISIM_NET_43),
                .Input_3(s_LOGISIM_NET_245),
                .Input_4(s_LOGISIM_NET_266),
                .Input_5(s_LOGISIM_NET_173),
                .Input_6(s_LOGISIM_NET_9),
                .Input_7(s_LOGISIM_NET_37),
                .Input_8(s_LOGISIM_NET_259),
                .Result(s_LOGISIM_NET_239));

   NOT_GATE      GATE_379 (.Input_1(s_LOGISIM_NET_7),
                           .Result(s_LOGISIM_NET_364));

   NOT_GATE      GATE_380 (.Input_1(s_LOGISIM_NET_31),
                           .Result(s_LOGISIM_NET_115));

   NOT_GATE      GATE_381 (.Input_1(s_LOGISIM_NET_32),
                           .Result(s_LOGISIM_NET_357));

   NOT_GATE      GATE_382 (.Input_1(s_LOGISIM_NET_7),
                           .Result(s_LOGISIM_NET_351));

   NOT_GATE      GATE_383 (.Input_1(s_LOGISIM_NET_18),
                           .Result(s_LOGISIM_NET_67));

   NOT_GATE      GATE_384 (.Input_1(s_LOGISIM_NET_31),
                           .Result(s_LOGISIM_NET_113));

   NOT_GATE      GATE_385 (.Input_1(s_LOGISIM_NET_14),
                           .Result(s_LOGISIM_NET_195));

   NOT_GATE      GATE_386 (.Input_1(s_LOGISIM_NET_10),
                           .Result(s_LOGISIM_NET_244));

   AND_GATE_8_INPUTS #(.BubblesMask(0))
      GATE_387 (.Input_1(s_LOGISIM_NET_187),
                .Input_2(s_LOGISIM_NET_0),
                .Input_3(s_LOGISIM_NET_9),
                .Input_4(s_LOGISIM_NET_32),
                .Input_5(s_LOGISIM_NET_210),
                .Input_6(s_LOGISIM_NET_7),
                .Input_7(s_LOGISIM_NET_263),
                .Input_8(s_LOGISIM_NET_75),
                .Result(s_LOGISIM_NET_251));

   NOT_GATE      GATE_388 (.Input_1(s_LOGISIM_NET_22),
                           .Result(s_LOGISIM_NET_0));

   AND_GATE_8_INPUTS #(.BubblesMask(0))
      GATE_389 (.Input_1(s_LOGISIM_NET_90),
                .Input_2(s_LOGISIM_NET_16),
                .Input_3(s_LOGISIM_NET_9),
                .Input_4(s_LOGISIM_NET_390),
                .Input_5(s_LOGISIM_NET_223),
                .Input_6(s_LOGISIM_NET_68),
                .Input_7(s_LOGISIM_NET_225),
                .Input_8(s_LOGISIM_NET_352),
                .Result(s_LOGISIM_NET_204));

   AND_GATE_8_INPUTS #(.BubblesMask(0))
      GATE_390 (.Input_1(s_LOGISIM_NET_5),
                .Input_2(s_LOGISIM_NET_7),
                .Input_3(s_LOGISIM_NET_321),
                .Input_4(s_LOGISIM_NET_403),
                .Input_5(s_LOGISIM_NET_324),
                .Input_6(s_LOGISIM_NET_9),
                .Input_7(s_LOGISIM_NET_253),
                .Input_8(s_LOGISIM_NET_110),
                .Result(s_LOGISIM_NET_112));

   NOT_GATE      GATE_391 (.Input_1(s_LOGISIM_NET_22),
                           .Result(s_LOGISIM_NET_339));

   AND_GATE_10_INPUTS #(.BubblesMask(0))
      GATE_392 (.Input_1(s_LOGISIM_NET_18),
                .Input_10(s_LOGISIM_NET_19),
                .Input_2(s_LOGISIM_NET_129),
                .Input_3(s_LOGISIM_NET_347),
                .Input_4(s_LOGISIM_NET_233),
                .Input_5(s_LOGISIM_NET_260),
                .Input_6(s_LOGISIM_NET_98),
                .Input_7(s_LOGISIM_NET_32),
                .Input_8(s_LOGISIM_NET_9),
                .Input_9(s_LOGISIM_NET_196),
                .Result(s_LOGISIM_NET_85));

   NOT_GATE      GATE_393 (.Input_1(s_LOGISIM_NET_35),
                           .Result(s_LOGISIM_NET_228));

   AND_GATE_8_INPUTS #(.BubblesMask(0))
      GATE_394 (.Input_1(s_LOGISIM_NET_76),
                .Input_2(s_LOGISIM_NET_272),
                .Input_3(s_LOGISIM_NET_107),
                .Input_4(s_LOGISIM_NET_32),
                .Input_5(s_LOGISIM_NET_378),
                .Input_6(s_LOGISIM_NET_344),
                .Input_7(s_LOGISIM_NET_7),
                .Input_8(s_LOGISIM_NET_118),
                .Result(s_LOGISIM_NET_386));



endmodule
